* NGSPICE file created from user_project_wrapper.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_4 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_4 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

.subckt user_project_wrapper io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
X_1270_ mprj.PS_Rx_inst6.LUT_inst1.i3 _0600_ _1270_/VDD _1270_/VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_1399_ _0014_ net71 mprj.PS_R1_inst1.LUT_inst14.I1 _1399_/VDD _1399_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0985_ _0296_ _0299_ _0327_ _0328_ net40 _0985_/VDD _0985_/VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_1184_ _0297_ _0204_ _0222_ _0269_ _0518_ _0519_ _1184_/VDD _1184_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0968_ _0279_ _0309_ _0311_ _0312_ _0968_/VDD _0968_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_4
X_1253_ _0249_ _0583_ _0584_ _1253_/VDD _1253_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0770_ _0104_ _0121_ _0122_ _0770_/VDD _0770_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1322_ _0641_ _0003_ _1322_/VDD _1322_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0899_ _0187_ mprj.PS_Rx_inst6.LUT_inst1.i3 _0245_ _0899_/VDD _0899_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_0753_ _0104_ _0068_ _0105_ _0753_/VDD _0753_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0822_ net8 _0170_ _0040_ _0171_ _0822_/VDD _0822_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0684_ net7 _0041_ _0684_/VDD _0684_/VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1305_ _0322_ mprj.PS_Rx_inst8.LUT_inst1.i3 _0631_ _1305_/VDD _1305_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1098_ _0147_ _0249_ _0289_ _0437_ _1098_/VDD _1098_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1167_ _0136_ mprj.PS_Rx_inst3.LUT_inst1.i3 _0451_ _0503_ _1167_/VDD _1167_/VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1236_ _0270_ _0323_ _0334_ _0568_ _1236_/VDD _1236_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1219_ _0190_ _0382_ _0443_ _0170_ _0551_ _0552_ _1219_/VDD _1219_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1021_ _0239_ _0116_ _0132_ _0216_ _0362_ _0363_ _1021_/VDD _1021_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0736_ _0067_ _0089_ _0050_ _0090_ _0736_/VDD _0736_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0805_ _0104_ mprj.PS_Rx_inst4.LUT_inst1.i3 _0155_ _0805_/VDD _0805_/VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
Xuser_project_wrapper_92 io_oeb[20] user_project_wrapper_92/VDD user_project_wrapper_92/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1004_ mprj.PS_R1_inst1.LUT_inst10.I1 _0119_ _0129_ _0347_ _1004_/VDD _1004_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xuser_project_wrapper_81 io_oeb[9] user_project_wrapper_81/VDD user_project_wrapper_81/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0719_ _0046_ _0065_ _0073_ _0719_/VDD _0719_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xuser_project_wrapper_119 io_out[12] user_project_wrapper_119/VDD user_project_wrapper_119/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xoutput53 net53 wbs_dat_o[25] output53/VDD output53/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput42 net42 wbs_dat_o[15] output42/VDD output42/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput64 net64 wbs_dat_o[6] output64/VDD output64/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xuser_project_wrapper_108 io_oeb[36] user_project_wrapper_108/VDD user_project_wrapper_108/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1398_ _0013_ net68 mprj.PS_R1_inst1.LUT_inst13.I1 _1398_/VDD _1398_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0984_ _0315_ _0326_ _0102_ _0328_ _0984_/VDD _1263_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1252_ _0237_ _0390_ _0244_ _0583_ _1252_/VDD _1252_/VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1321_ net23 _0071_ _0637_ _0641_ _1321_/VDD _1321_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1183_ _0297_ _0209_ _0220_ _0518_ _1183_/VDD _1183_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0967_ mprj.PS_R1_inst1.LUT_inst11.I1 _0076_ _0138_ mprj.PS_R1_inst1.LUT_inst10.I1
+ _0310_ _0311_ _0967_/VDD _0967_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0898_ _0187_ mprj.PS_Rx_inst6.LUT_inst1.i3 _0244_ _0898_/VDD _0898_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0821_ _0169_ _0170_ _0821_/VDD _0821_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_0752_ mprj.PS_Rx_inst3.LUT_inst1.i4 _0104_ _0752_/VDD _0752_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1097_ _0433_ _0435_ _0436_ _1097_/VDD _1097_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1304_ _0630_ net57 _1304_/VDD _1304_/VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1235_ _0217_ _0382_ _0443_ _0190_ _0566_ _0567_ _1235_/VDD _1235_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0683_ _0036_ _0038_ _0039_ _0040_ _0683_/VDD _0683_/VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_1166_ _0486_ _0501_ _0502_ _1166_/VDD _1166_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_1020_ mprj.PS_R1_inst1.LUT_inst11.I1 _0119_ _0130_ _0362_ _1020_/VDD _1020_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0804_ mprj.PS_Rx_inst4.LUT_inst1.i4 _0154_ _0804_/VDD _0804_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_0735_ _0085_ _0088_ _0089_ _0735_/VDD _0735_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1149_ _0086_ _0454_ _0485_ _0486_ _1149_/VDD _1149_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1218_ _0190_ _0385_ _0411_ _0551_ _1218_/VDD _1218_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xuser_project_wrapper_93 io_oeb[21] user_project_wrapper_93/VDD user_project_wrapper_93/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1003_ _0169_ _0156_ _0175_ _0146_ _0345_ _0346_ _1003_/VDD _1003_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xuser_project_wrapper_82 io_oeb[10] user_project_wrapper_82/VDD user_project_wrapper_82/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0718_ _0058_ _0071_ _0064_ _0072_ _0718_/VDD _0718_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xoutput54 net54 wbs_dat_o[26] output54/VDD output54/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput43 net43 wbs_dat_o[16] output43/VDD output43/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput65 net65 wbs_dat_o[7] output65/VDD output65/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xuser_project_wrapper_109 io_oeb[37] user_project_wrapper_109/VDD user_project_wrapper_109/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xoutput32 net32 io_out[0] output32/VDD output32/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_0983_ _0315_ _0326_ _0327_ _0983_/VDD _0983_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
X_1397_ _0012_ net71 mprj.PS_R1_inst1.LUT_inst12.I1 _1397_/VDD _1397_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_1320_ _0640_ _0002_ _1320_/VDD _1320_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1182_ _0147_ _0382_ _0443_ _0127_ _0516_ _0517_ _1182_/VDD _1182_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1251_ _0298_ _0320_ _0337_ _0270_ _0581_ _0582_ _1251_/VDD _1251_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0897_ mprj.PS_Rx_inst6.LUT_inst1.i3 _0237_ _0243_ _0897_/VDD _0897_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_0966_ mprj.PS_R1_inst1.LUT_inst11.I1 _0081_ _0099_ _0310_ _0966_/VDD _0966_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1234_ _0217_ _0385_ _0411_ _0566_ _1234_/VDD _1234_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1165_ _0330_ _0157_ _0175_ _0297_ _0500_ _0501_ _1165_/VDD _1165_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0682_ net7 _0032_ _0039_ _0682_/VDD _0682_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1303_ _0627_ _0628_ _0629_ _0630_ _1303_/VDD _1303_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1096_ _0189_ _0205_ _0222_ _0169_ _0434_ _0435_ _1096_/VDD _1096_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0751_ _0092_ _0095_ _0101_ _0103_ net62 _0751_/VDD _0751_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_0820_ mprj.PS_R1_inst1.LUT_inst8.I1 _0169_ _0820_/VDD _0820_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0949_ _0282_ _0292_ _0293_ _0294_ _0949_/VDD _0949_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0803_ _0078_ _0104_ _0149_ _0150_ _0152_ _0153_ _0803_/VDD _0803_/VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_0734_ _0086_ _0077_ _0087_ _0088_ _0734_/VDD _0734_/VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_1079_ _0377_ _0417_ _0103_ _0419_ _1079_/VDD _1079_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1148_ _0449_ _0116_ _0132_ _0483_ _0484_ _0485_ _1148_/VDD _1148_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1217_ _0051_ _0550_ net50 _1217_/VDD _1217_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xuser_project_wrapper_94 io_oeb[22] user_project_wrapper_94/VDD user_project_wrapper_94/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0717_ _0070_ _0071_ _0717_/VDD _0717_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
Xuser_project_wrapper_83 io_oeb[11] user_project_wrapper_83/VDD user_project_wrapper_83/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1002_ _0169_ _0152_ _0173_ _0345_ _1002_/VDD _1002_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xuser_project_wrapper_72 io_oeb[0] user_project_wrapper_72/VDD user_project_wrapper_72/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xoutput55 net55 wbs_dat_o[27] output55/VDD output55/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput44 net44 wbs_dat_o[17] output44/VDD output44/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput66 net66 wbs_dat_o[8] output66/VDD output66/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net33 io_out[1] output33/VDD output33/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_0982_ _0295_ _0325_ _0326_ _0982_/VDD _0982_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_1396_ _0011_ net71 mprj.PS_R1_inst1.LUT_inst11.I1 _1396_/VDD _1396_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0965_ _0189_ _0115_ _0131_ _0169_ _0308_ _0309_ _0965_/VDD _0965_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1181_ _0147_ _0385_ _0411_ _0516_ _1181_/VDD _1181_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0896_ mprj.PS_Rx_inst6.LUT_inst1.i4 _0242_ _0896_/VDD _0896_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_1250_ _0298_ _0323_ _0334_ _0581_ _1250_/VDD _1250_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1379_ net19 mprj.PS_Rx_inst8.LUT_inst1.i3 _0655_ _0672_ _1379_/VDD _1379_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1302_ _0627_ _0628_ _0051_ _0629_ _1302_/VDD _1302_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0681_ net31 _0037_ _0038_ _0681_/VDD _0681_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1233_ _0421_ _0565_ net51 _1233_/VDD _1233_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1095_ _0189_ _0209_ _0220_ _0434_ _1095_/VDD _1095_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1164_ _0330_ _0152_ _0173_ _0500_ _1164_/VDD _1164_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0750_ _0102_ _0103_ _0750_/VDD _0750_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_0948_ _0282_ _0292_ _0050_ _0293_ _0948_/VDD _0948_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0879_ _0126_ _0119_ _0130_ _0226_ _0879_/VDD _0879_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0802_ _0151_ _0152_ _0802_/VDD _0802_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0733_ _0052_ _0065_ _0067_ _0078_ _0087_ _0733_/VDD _0733_/VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_1078_ _0377_ _0417_ _0418_ _1078_/VDD _1078_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1216_ _0530_ _0547_ _0549_ _0550_ _1216_/VDD _1216_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1147_ _0449_ _0130_ _0484_ _1147_/VDD _1147_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0716_ mprj.PS_R1_inst1.LUT_inst3.I1 _0070_ _0716_/VDD _0716_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
Xuser_project_wrapper_95 io_oeb[23] user_project_wrapper_95/VDD user_project_wrapper_95/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_84 io_oeb[12] user_project_wrapper_84/VDD user_project_wrapper_84/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1001_ _0126_ _0204_ _0221_ mprj.PS_R1_inst1.LUT_inst5.I1 _0343_ _0344_ _1001_/VDD
+ _1001_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xuser_project_wrapper_73 io_oeb[1] user_project_wrapper_73/VDD user_project_wrapper_73/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xoutput56 net56 wbs_dat_o[28] output56/VDD output56/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput45 net45 wbs_dat_o[18] output45/VDD output45/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput67 net67 wbs_dat_o[9] output67/VDD output67/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[2] output34/VDD output34/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_0981_ _0059_ _0320_ _0321_ _0250_ _0324_ _0325_ _0981_/VDD _0981_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1395_ _0010_ net69 mprj.PS_R1_inst1.LUT_inst10.I1 _1395_/VDD _1395_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_1180_ _0051_ _0515_ net48 _1180_/VDD _1180_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0895_ _0058_ _0240_ _0064_ _0241_ _0895_/VDD _0895_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0964_ mprj.PS_R1_inst1.LUT_inst10.I0 _0119_ _0129_ _0308_ _0964_/VDD _0964_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1378_ _0322_ _0656_ _0671_ _0029_ _1378_/VDD _1378_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1301_ _0086_ _0620_ _0628_ _1301_/VDD _1301_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_0680_ net13 net30 _0037_ _0680_/VDD _0680_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1232_ _0547_ _0563_ _0564_ _0565_ _1232_/VDD _1232_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0947_ _0265_ _0291_ _0292_ _0947_/VDD _0947_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_1094_ _0403_ _0430_ _0432_ _0433_ _1094_/VDD _1094_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_1163_ _0217_ _0247_ _0286_ _0190_ _0498_ _0499_ _1163_/VDD _1163_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_0878_ _0063_ _0220_ _0223_ _0224_ _0225_ _0878_/VDD _0878_/VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1077_ _0409_ _0416_ _0417_ _1077_/VDD _1077_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_1215_ _0170_ _0382_ _0443_ _0147_ _0548_ _0549_ _1215_/VDD _1215_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1146_ mprj.PS_R1_inst1.LUT_inst14.I1 _0117_ _0483_ _1146_/VDD _1146_/VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
X_0801_ _0104_ mprj.PS_Rx_inst4.LUT_inst1.i3 _0151_ _0801_/VDD _0801_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_0732_ _0046_ _0048_ _0086_ _0732_/VDD _0732_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_project_wrapper_96 io_oeb[24] user_project_wrapper_96/VDD user_project_wrapper_96/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_85 io_oeb[13] user_project_wrapper_85/VDD user_project_wrapper_85/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0715_ _0067_ _0068_ _0069_ _0715_/VDD _0715_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1000_ _0126_ _0208_ _0219_ _0343_ _1000_/VDD _1000_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xuser_project_wrapper_74 io_oeb[2] user_project_wrapper_74/VDD user_project_wrapper_74/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1129_ _0436_ _0463_ _0466_ _0467_ _1129_/VDD _1129_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
Xoutput57 net57 wbs_dat_o[29] output57/VDD output57/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput46 net46 wbs_dat_o[19] output46/VDD output46/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 wbs_ack_o output35/VDD output35/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_0980_ _0035_ _0322_ _0323_ _0324_ _0980_/VDD _0980_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1394_ _0009_ net69 mprj.PS_R1_inst1.LUT_inst10.I0 _1394_/VDD _1394_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0963_ _0146_ _0156_ _0174_ mprj.PS_R1_inst1.LUT_inst6.I1 _0306_ _0307_ _0963_/VDD
+ _0963_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0894_ _0239_ _0240_ _0894_/VDD _0894_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1377_ net18 _0657_ _0671_ _1377_/VDD _1377_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xfanout70 net71 net70 fanout70/VDD _1407_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_0946_ _0062_ _0248_ _0284_ _0287_ _0290_ _0291_ _0946_/VDD _0946_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1231_ _0547_ _0563_ _0051_ _0564_ _1231_/VDD _1231_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1093_ _0239_ _0157_ _0175_ _0216_ _0431_ _0432_ _1093_/VDD _1093_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1300_ _0586_ _0411_ _0625_ _0626_ _0627_ _1300_/VDD _1300_/VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1162_ _0216_ _0249_ _0288_ _0498_ _1162_/VDD _1162_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0877_ _0063_ _0205_ _0224_ _0877_/VDD _0877_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1214_ _0170_ _0385_ _0411_ _0548_ _1214_/VDD _1214_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1145_ _0426_ _0481_ _0482_ _1145_/VDD _1145_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_0731_ _0084_ _0085_ _0731_/VDD _0731_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_0800_ _0078_ _0144_ _0150_ _0800_/VDD _0800_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_0929_ mprj.PS_R1_inst1.LUT_inst6.I1 _0152_ _0172_ _0274_ _0929_/VDD _0929_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1076_ _0062_ _0411_ _0414_ _0415_ _0416_ _1076_/VDD _1076_/VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xuser_project_wrapper_86 io_oeb[14] user_project_wrapper_86/VDD user_project_wrapper_86/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_97 io_oeb[25] user_project_wrapper_97/VDD user_project_wrapper_97/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_75 io_oeb[3] user_project_wrapper_75/VDD user_project_wrapper_75/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1128_ _0404_ _0465_ _0466_ _1128_/VDD _1128_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1059_ mprj.PS_R1_inst1.LUT_inst12.I1 _0119_ _0130_ _0399_ _1059_/VDD _1059_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0714_ _0043_ _0068_ _0714_/VDD _0714_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
Xoutput58 net58 wbs_dat_o[2] output58/VDD output58/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput47 net47 wbs_dat_o[1] output47/VDD output47/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput36 net36 wbs_dat_o[0] output36/VDD output36/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1393_ _0008_ net69 mprj.PS_R1_inst1.LUT_inst8.I1 _1393_/VDD _1393_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0893_ mprj.PS_R1_inst1.LUT_inst11.I1 _0239_ _0893_/VDD _0893_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1376_ _0373_ _0656_ _0670_ _0028_ _1376_/VDD _1376_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0962_ _0146_ _0151_ _0172_ _0306_ _0962_/VDD _0962_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xfanout71 net3 net71 _1399_/VDD fanout71/VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_1092_ _0239_ _0152_ _0173_ _0431_ _1092_/VDD _1092_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1230_ _0552_ _0562_ _0563_ _1230_/VDD _1230_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_0876_ _0059_ _0206_ _0222_ _0223_ _0876_/VDD _0876_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1161_ _0170_ _0319_ _0337_ _0147_ _0496_ _0497_ _1161_/VDD _1161_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0945_ _0062_ _0289_ _0290_ _0945_/VDD _0945_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1359_ net24 mprj.PS_Rx_inst3.LUT_inst1.i3 _0655_ _0662_ _1359_/VDD _1359_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1213_ _0527_ _0535_ _0546_ _0547_ _1213_/VDD _1213_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_4
X_0730_ _0046_ _0054_ _0077_ _0083_ _0084_ _0730_/VDD _0730_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_1144_ _0297_ _0156_ _0174_ _0269_ _0480_ _0481_ _1144_/VDD _1144_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0859_ mprj.PS_R1_inst1.LUT_inst1.i0 _0187_ _0207_ _0859_/VDD _0859_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0928_ _0093_ _0205_ _0222_ mprj.PS_R1_inst1.LUT_inst3.I1 _0272_ _0273_ _0928_/VDD
+ _0928_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1075_ _0062_ _0381_ _0415_ _1075_/VDD _1075_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xuser_project_wrapper_87 io_oeb[15] user_project_wrapper_87/VDD user_project_wrapper_87/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_98 io_oeb[26] user_project_wrapper_98/VDD user_project_wrapper_98/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_76 io_oeb[4] user_project_wrapper_76/VDD user_project_wrapper_76/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1127_ _0170_ _0247_ _0286_ _0146_ _0464_ _0465_ _1127_/VDD _1127_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1058_ _0216_ _0157_ _0175_ _0189_ _0397_ _0398_ _1058_/VDD _1058_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0713_ mprj.PS_Rx_inst2.LUT_inst1.i4 _0067_ _0713_/VDD _0713_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
Xoutput59 net59 wbs_dat_o[30] output59/VDD output59/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput48 net48 wbs_dat_o[20] output48/VDD output48/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput37 net37 wbs_dat_o[10] output37/VDD output37/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1392_ _0007_ net68 mprj.PS_R1_inst1.LUT_inst7.I1 _1392_/VDD _1392_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0892_ _0237_ _0068_ _0238_ _0892_/VDD _0892_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1375_ net17 _0657_ _0670_ _1375_/VDD _1375_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0961_ _0106_ _0204_ _0221_ mprj.PS_R1_inst1.LUT_inst4.I1 _0304_ _0305_ _0961_/VDD
+ _0961_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0944_ _0288_ _0289_ _0944_/VDD _0944_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1160_ _0170_ _0323_ _0333_ _0496_ _1160_/VDD _1160_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1091_ _0426_ _0429_ _0430_ _1091_/VDD _1091_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_0875_ _0221_ _0222_ _0875_/VDD _0875_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1358_ _0136_ _0656_ _0661_ _0019_ _1358_/VDD _1358_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1289_ _0331_ _0381_ _0413_ _0298_ _0616_ _0617_ _1289_/VDD _1289_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0927_ _0093_ _0209_ _0220_ _0272_ _0927_/VDD _0927_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1074_ mprj.PS_R1_inst1.LUT_inst1.i1 _0383_ _0413_ _0414_ _1074_/VDD _1074_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0858_ mprj.PS_Rx_inst5.LUT_inst1.i3 _0187_ _0206_ _0858_/VDD _0858_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_1212_ _0524_ _0537_ _0545_ _0546_ _1212_/VDD _1212_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1143_ _0297_ _0151_ _0172_ _0480_ _1143_/VDD _1143_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0789_ _0094_ _0076_ _0138_ _0070_ _0139_ _0140_ _0789_/VDD _0789_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xuser_project_wrapper_88 io_oeb[16] user_project_wrapper_88/VDD user_project_wrapper_88/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_99 io_oeb[27] user_project_wrapper_99/VDD user_project_wrapper_99/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0712_ _0052_ _0048_ _0051_ _0066_ net58 _0712_/VDD _0712_/VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
Xuser_project_wrapper_77 io_oeb[5] user_project_wrapper_77/VDD user_project_wrapper_77/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1126_ _0169_ _0245_ _0288_ _0464_ _1126_/VDD _1126_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1057_ _0216_ _0152_ _0173_ _0397_ _1057_/VDD _1057_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xoutput49 net49 wbs_dat_o[21] output49/VDD output49/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput38 net38 wbs_dat_o[11] output38/VDD output38/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1109_ _0127_ _0323_ _0334_ _0447_ _1109_/VDD _1109_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1391_ _0006_ net68 mprj.PS_R1_inst1.LUT_inst6.I1 _1391_/VDD _1391_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0891_ mprj.PS_Rx_inst6.LUT_inst1.i4 _0237_ _0891_/VDD _0891_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
Xuser_project_wrapper_210 user_irq[1] user_project_wrapper_210/VDD user_project_wrapper_210/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0960_ mprj.PS_R1_inst1.LUT_inst5.I1 _0209_ _0219_ _0304_ _0960_/VDD _0960_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1374_ _0242_ _0656_ _0669_ _0027_ _1374_/VDD _1374_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1090_ _0402_ _0428_ _0429_ _1090_/VDD _1090_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1357_ net23 _0657_ _0661_ _1357_/VDD _1357_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0874_ _0201_ _0202_ _0208_ _0221_ _0874_/VDD _0874_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0943_ _0187_ mprj.PS_Rx_inst6.LUT_inst1.i3 mprj.PS_Rx_inst6.LUT_inst1.i4 _0288_
+ _0943_/VDD _0943_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1288_ _0331_ _0378_ _0410_ _0616_ _1288_/VDD _1288_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1142_ _0190_ _0248_ _0287_ _0170_ _0478_ _0479_ _1142_/VDD _1142_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0926_ _0058_ _0270_ _0064_ _0271_ _0926_/VDD _0926_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1211_ _0523_ _0544_ _0545_ _1211_/VDD _1211_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1073_ _0378_ _0412_ _0413_ _1073_/VDD _1073_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_0857_ _0204_ _0205_ _0857_/VDD _0857_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1409_ _0024_ net70 mprj.PS_Rx_inst5.LUT_inst1.i3 _1409_/VDD _1409_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0788_ _0094_ _0081_ _0099_ _0139_ _0788_/VDD _0788_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xuser_project_wrapper_89 io_oeb[17] user_project_wrapper_89/VDD user_project_wrapper_89/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_78 io_oeb[6] user_project_wrapper_78/VDD user_project_wrapper_78/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0711_ _0063_ _0064_ _0043_ _0065_ _0051_ _0066_ _0711_/VDD _0711_/VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_1056_ _0127_ _0248_ _0287_ _0107_ _0395_ _0396_ _1056_/VDD _1056_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0909_ _0106_ _0157_ _0175_ mprj.PS_R1_inst1.LUT_inst4.I1 _0254_ _0255_ _0909_/VDD
+ _0909_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xoutput39 net39 wbs_dat_o[12] output39/VDD output39/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1125_ _0433_ _0460_ _0462_ _0463_ _1125_/VDD _1125_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1039_ _0378_ _0380_ _0381_ _1039_/VDD _1039_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_1108_ _0051_ _0446_ net44 _1108_/VDD _1108_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1390_ _0005_ net70 mprj.PS_R1_inst1.LUT_inst5.I1 _1390_/VDD _1390_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0890_ _0215_ _0218_ _0235_ _0236_ net37 _0890_/VDD _0890_/VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
Xuser_project_wrapper_200 la_data_out[55] user_project_wrapper_200/VDD user_project_wrapper_200/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_211 user_irq[2] user_project_wrapper_211/VDD user_project_wrapper_211/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1373_ net16 _0657_ _0669_ _1373_/VDD _1373_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_0942_ _0286_ _0287_ _0974_/VDD _0942_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0873_ _0219_ _0220_ _0873_/VDD _0873_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1356_ _0660_ _0018_ _1356_/VDD _1356_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1287_ _0421_ _0615_ net55 _1287_/VDD _1287_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1072_ mprj.PS_Rx_inst8.LUT_inst1.i4 _0379_ _0412_ _1072_/VDD _1072_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1210_ _0506_ _0539_ _0543_ _0544_ _1210_/VDD _1210_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1141_ _0189_ _0249_ _0289_ _0478_ _1141_/VDD _1141_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0856_ _0144_ mprj.PS_Rx_inst5.LUT_inst1.i3 _0203_ _0204_ _0856_/VDD _0856_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1408_ _0023_ net70 mprj.PS_Rx_inst4.LUT_inst1.i4 _1408_/VDD _1408_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0787_ _0137_ _0138_ _0787_/VDD _0787_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0925_ _0269_ _0270_ _0925_/VDD _0925_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1339_ _0650_ _0011_ _1339_/VDD _1339_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xuser_project_wrapper_79 io_oeb[7] user_project_wrapper_79/VDD user_project_wrapper_79/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0710_ mprj.PS_Rx_inst2.LUT_inst1.i3 _0065_ _0710_/VDD _0710_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1055_ _0126_ _0249_ _0289_ _0395_ _1055_/VDD _1055_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1124_ _0216_ _0205_ _0222_ _0189_ _0461_ _0462_ _1124_/VDD _1124_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0839_ mprj.PS_Rx_inst5.LUT_inst1.i4 _0187_ _0839_/VDD _0839_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0908_ _0106_ _0152_ _0173_ _0254_ _0908_/VDD _0908_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1038_ mprj.PS_Rx_inst8.LUT_inst1.i4 _0379_ _0380_ _1038_/VDD _1038_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1107_ _0409_ _0441_ _0445_ _0446_ _1107_/VDD _1107_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1372_ _0600_ _0656_ _0668_ _0026_ _1372_/VDD _1372_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xuser_project_wrapper_201 la_data_out[56] user_project_wrapper_201/VDD user_project_wrapper_201/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1355_ net22 _0065_ _0655_ _0660_ _1355_/VDD _1355_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0941_ _0245_ _0285_ _0286_ _0941_/VDD _0941_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_0872_ _0187_ _0202_ _0219_ _0872_/VDD _0872_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1286_ _0597_ _0613_ _0614_ _0615_ _1286_/VDD _1286_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1140_ _0147_ _0320_ _0337_ _0127_ _0476_ _0477_ _1140_/VDD _1140_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1071_ _0410_ _0411_ _1071_/VDD _1071_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1269_ _0270_ _0381_ _0413_ _0240_ _0598_ _0599_ _1269_/VDD _1269_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1338_ net16 _0240_ _0642_ _0650_ _1338_/VDD _1338_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1407_ _0022_ net70 mprj.PS_Rx_inst4.LUT_inst1.i3 _1407_/VDD _1407_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0786_ _0136_ _0079_ _0080_ _0137_ _0786_/VDD _0786_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0855_ _0201_ _0202_ _0203_ _0855_/VDD _0855_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_0924_ mprj.PS_R1_inst1.LUT_inst12.I1 _0269_ _0924_/VDD _0924_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1123_ _0216_ _0209_ _0220_ _0461_ _1123_/VDD _1123_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1054_ _0094_ _0319_ _0336_ _0070_ _0393_ _0394_ _1054_/VDD _1054_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0907_ _0242_ _0252_ _0253_ _0907_/VDD _0907_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_0838_ _0168_ _0171_ _0186_ net66 _0838_/VDD _0838_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0769_ _0059_ _0116_ _0120_ _0121_ _0769_/VDD _0769_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1106_ _0071_ _0411_ _0442_ _0444_ _0445_ _1106_/VDD _1106_/VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1037_ _0295_ mprj.PS_Rx_inst8.LUT_inst1.i3 _0379_ _1037_/VDD _1037_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1371_ net15 _0657_ _0668_ _1371_/VDD _1371_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xuser_project_wrapper_202 la_data_out[57] user_project_wrapper_202/VDD user_project_wrapper_202/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0871_ _0058_ _0217_ _0064_ _0218_ _0871_/VDD _0871_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0940_ mprj.PS_Rx_inst6.LUT_inst1.i4 _0244_ _0285_ _0940_/VDD _0940_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1354_ _0052_ _0656_ _0659_ _0017_ _1354_/VDD _1354_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1285_ _0597_ _0613_ _0050_ _0614_ _1285_/VDD _1285_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1406_ _0021_ net70 mprj.PS_Rx_inst3.LUT_inst1.i4 _1406_/VDD _1406_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1070_ _0295_ mprj.PS_Rx_inst8.LUT_inst1.i3 mprj.PS_Rx_inst8.LUT_inst1.i4 _0410_
+ _1070_/VDD _1070_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1337_ _0649_ _0010_ _1337_/VDD _1337_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0854_ mprj.PS_Rx_inst4.LUT_inst1.i4 mprj.PS_Rx_inst5.LUT_inst1.i3 _0202_ _0854_/VDD
+ _0854_/VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
X_0923_ mprj.PS_Rx_inst7.LUT_inst1.i3 _0068_ _0268_ _0923_/VDD _0923_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0785_ mprj.PS_Rx_inst2.LUT_inst1.i4 _0136_ _0785_/VDD _0785_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_1268_ _0270_ _0378_ _0410_ _0598_ _1268_/VDD _1268_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1199_ _0051_ _0532_ _0533_ _0420_ net49 _1199_/VDD _1199_/VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_1053_ _0094_ _0316_ _0333_ _0393_ _1053_/VDD _1053_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1122_ _0429_ _0457_ _0459_ _0460_ _1122_/VDD _1122_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_0837_ _0178_ _0184_ _0185_ _0186_ _0837_/VDD _0837_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0768_ _0078_ _0067_ _0117_ _0118_ _0119_ _0120_ _0768_/VDD _0768_/VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_0699_ _0052_ _0054_ _0055_ _0699_/VDD _0699_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0906_ _0207_ _0243_ _0248_ _0059_ _0251_ _0252_ _0906_/VDD _0906_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1105_ _0062_ _0383_ _0443_ _0444_ _1105_/VDD _1105_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1036_ _0295_ mprj.PS_Rx_inst8.LUT_inst1.i3 _0378_ _1036_/VDD _1036_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1019_ _0189_ _0156_ _0174_ _0169_ _0360_ _0361_ _1019_/VDD _1019_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1370_ _0201_ _0656_ _0667_ _0025_ _1370_/VDD _1370_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xuser_project_wrapper_203 la_data_out[58] user_project_wrapper_203/VDD user_project_wrapper_203/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0870_ _0216_ _0217_ _0870_/VDD _0870_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1284_ _0608_ _0612_ _0613_ _1284_/VDD _1284_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_0999_ _0093_ _0247_ _0286_ mprj.PS_R1_inst1.LUT_inst3.I1 _0341_ _0342_ _0999_/VDD
+ _0999_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1353_ net21 _0657_ _0659_ _1353_/VDD _1353_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0853_ _0187_ _0201_ _0853_/VDD _0853_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_1405_ _0020_ net68 mprj.PS_Rx_inst3.LUT_inst1.i3 _1405_/VDD _1405_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0922_ _0238_ _0241_ _0266_ _0267_ net38 _0922_/VDD _0922_/VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_0784_ _0063_ _0130_ _0133_ _0134_ _0135_ _0784_/VDD _0784_/VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1198_ _0512_ _0531_ _0533_ _1198_/VDD _1198_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
X_1267_ _0590_ _0596_ _0597_ _1267_/VDD _1267_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
Xinput1 io_in[2] net1 input1/VDD input1/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1336_ net15 _0217_ _0642_ _0649_ _1336_/VDD _1336_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1121_ _0269_ _0157_ _0175_ _0239_ _0458_ _0459_ _1121_/VDD _1121_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1052_ _0389_ _0392_ net42 _1052_/VDD _1052_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0767_ _0113_ _0119_ _0767_/VDD _0999_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0905_ _0249_ _0250_ _0251_ _0905_/VDD _0905_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1319_ net22 _0063_ _0637_ _0640_ _1319_/VDD _1319_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0836_ _0178_ _0184_ _0102_ _0185_ _0836_/VDD _0836_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0698_ mprj.PS_R1_inst1.LUT_inst1.i0 _0053_ mprj.PS_R1_inst1.LUT_inst1.i3 _0054_
+ _0698_/VDD _0698_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1035_ _0354_ _0371_ _0376_ _0377_ _1035_/VDD _1035_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1104_ _0413_ _0443_ _1104_/VDD _1104_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0819_ mprj.PS_Rx_inst5.LUT_inst1.i3 _0044_ _0168_ _0819_/VDD _0819_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1018_ _0189_ _0152_ _0172_ _0360_ _1018_/VDD _1018_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xuser_project_wrapper_204 la_data_out[59] user_project_wrapper_204/VDD user_project_wrapper_204/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1283_ _0055_ _0611_ _0612_ _1283_/VDD _1283_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_1352_ _0047_ _0656_ _0658_ _0016_ _1352_/VDD _1352_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0998_ mprj.PS_R1_inst1.LUT_inst4.I1 _0245_ _0288_ _0341_ _0998_/VDD _0998_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0921_ _0253_ _0265_ _0103_ _0267_ _0921_/VDD _0921_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0852_ _0183_ _0194_ _0199_ _0200_ _0852_/VDD _0852_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_0783_ _0063_ _0116_ _0134_ _0783_/VDD _0783_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1404_ _0019_ net69 mprj.PS_Rx_inst2.LUT_inst1.i4 _1404_/VDD _1404_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_1266_ _0331_ _0320_ _0337_ _0298_ _0595_ _0596_ _1266_/VDD _1266_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1197_ _0512_ _0531_ _0532_ _1197_/VDD _1197_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1335_ _0648_ _0009_ _1335_/VDD _1335_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput2 io_in[3] net2 input2/VDD input2/VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1318_ _0053_ _0637_ _0639_ _0001_ _1318_/VDD _1318_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0766_ _0078_ _0104_ _0118_ _0766_/VDD _0766_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_0697_ mprj.PS_R1_inst1.LUT_inst1.i1 _0053_ _0697_/VDD _0697_/VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_0835_ _0165_ _0183_ _0184_ _0835_/VDD _0835_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1051_ mprj.PS_Rx_inst8.LUT_inst1.i4 _0068_ _0391_ _0064_ _0392_ _1051_/VDD _1051_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_1120_ _0269_ _0152_ _0173_ _0458_ _1120_/VDD _1120_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0904_ _0078_ _0237_ _0250_ _0904_/VDD _0904_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1249_ _0240_ _0381_ _0443_ _0217_ _0579_ _0580_ _1249_/VDD _1249_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1034_ _0070_ _0334_ _0372_ _0375_ _0376_ _1034_/VDD _1034_/VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1103_ _0071_ _0382_ _0442_ _1103_/VDD _1103_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0749_ _0057_ _0060_ _0102_ _0749_/VDD _0749_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0818_ _0145_ _0148_ _0167_ net65 _0818_/VDD _0818_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1017_ _0106_ _0247_ _0286_ _0093_ _0358_ _0359_ _1017_/VDD _1017_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xuser_project_wrapper_205 la_data_out[60] user_project_wrapper_205/VDD user_project_wrapper_205/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xfanout68 net3 net68 fanout68/VDD _1410_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_1282_ _0586_ _0334_ _0609_ _0610_ _0611_ _1282_/VDD _1282_/VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1351_ net14 _0657_ _0658_ _1351_/VDD _1351_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_0997_ _0063_ _0334_ _0339_ _0340_ _0997_/VDD _0997_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0920_ _0253_ _0265_ _0266_ _0920_/VDD _0920_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_0851_ _0180_ _0196_ _0198_ _0199_ _0851_/VDD _0851_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_1196_ _0517_ _0530_ _0531_ _1196_/VDD _1196_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_1403_ _0018_ net69 mprj.PS_Rx_inst2.LUT_inst1.i3 _1403_/VDD _1403_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0782_ _0059_ _0117_ _0132_ _0133_ _0782_/VDD _0782_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1334_ net29 _0190_ _0642_ _0648_ _1334_/VDD _1334_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1265_ _0331_ _0323_ _0334_ _0595_ _1265_/VDD _1265_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xinput3 wb_clk_i net3 input3/VDD input3/VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_0834_ _0164_ _0180_ _0182_ _0183_ _0834_/VDD _0834_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_0765_ mprj.PS_Rx_inst3.LUT_inst1.i3 _0104_ _0117_ _0765_/VDD _0765_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_1050_ net8 _0390_ _0391_ _1050_/VDD _1050_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0696_ _0046_ _0052_ _0696_/VDD _0696_/VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
X_0903_ _0245_ _0249_ _0903_/VDD _0903_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1317_ net21 _0637_ _0639_ _1317_/VDD _1317_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1248_ _0240_ _0385_ _0410_ _0579_ _1248_/VDD _1248_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1179_ _0492_ _0512_ _0514_ _0515_ _1179_/VDD _1179_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1102_ _0408_ _0423_ _0440_ _0441_ _1102_/VDD _1102_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_0748_ _0063_ _0076_ _0100_ _0101_ _0748_/VDD _0748_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0817_ _0159_ _0165_ _0166_ _0167_ _0817_/VDD _0817_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1033_ mprj.PS_R1_inst1.LUT_inst2.I1 _0374_ _0336_ _0375_ _1033_/VDD _1033_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0679_ net6 net5 _0036_ _0679_/VDD _0679_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1016_ _0106_ _0245_ _0288_ _0358_ _1016_/VDD _1016_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xuser_project_wrapper_206 la_data_out[61] user_project_wrapper_206/VDD user_project_wrapper_206/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xfanout69 net3 net69 _1400_/VDD fanout69/VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1350_ _0655_ _0657_ _1350_/VDD _1350_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1281_ _0331_ _0374_ _0337_ _0610_ _1281_/VDD _1281_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0996_ _0062_ _0320_ _0337_ _0338_ _0339_ _0996_/VDD _0996_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_0781_ _0131_ _0132_ _0781_/VDD _0781_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1333_ _0647_ _0008_ _1333_/VDD _1333_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1264_ _0421_ _0594_ net53 _1264_/VDD _1264_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1402_ _0017_ net70 mprj.PS_R1_inst1.LUT_inst1.i4 _1402_/VDD _1402_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_1195_ _0511_ _0527_ _0529_ _0530_ _1195_/VDD _1195_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xinput4 wb_rst_i net4 input4/VDD input4/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_0850_ _0106_ _0116_ _0132_ mprj.PS_R1_inst1.LUT_inst4.I1 _0197_ _0198_ _1360_/VDD
+ _0850_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0979_ _0316_ _0323_ _0979_/VDD _0979_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0833_ _0093_ _0116_ _0132_ mprj.PS_R1_inst1.LUT_inst3.I1 _0181_ _0182_ _0833_/VDD
+ _0833_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0902_ _0247_ _0248_ _0902_/VDD _0902_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0695_ _0050_ _0051_ _0695_/VDD _0695_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1247_ _0562_ _0577_ _0578_ net52 _1247_/VDD _1247_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0764_ _0115_ _0116_ _0764_/VDD _0764_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1316_ _0035_ _0637_ _0638_ _0000_ _1316_/VDD _1316_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1178_ _0127_ _0382_ _0443_ _0107_ _0513_ _0514_ _1178_/VDD _1178_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0816_ _0159_ _0165_ _0050_ _0166_ _0816_/VDD _0816_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0678_ mprj.PS_R1_inst1.LUT_inst1.i0 _0035_ _0678_/VDD _0678_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_1032_ _0373_ _0322_ _0374_ _1032_/VDD _1032_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1101_ _0436_ _0439_ _0440_ _1101_/VDD _1101_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_0747_ _0096_ _0097_ _0099_ _0063_ _0100_ _0747_/VDD _0747_/VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_1015_ _0329_ _0332_ _0357_ net41 _1015_/VDD _1015_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xuser_project_wrapper_207 la_data_out[62] user_project_wrapper_207/VDD user_project_wrapper_207/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1280_ _0586_ _0320_ _0609_ _1280_/VDD _1280_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0995_ _0053_ _0321_ _0338_ _0995_/VDD _0995_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1194_ _0190_ _0320_ _0337_ _0170_ _0528_ _0529_ _1194_/VDD _1194_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0780_ _0112_ _0114_ _0113_ _0131_ _0780_/VDD _0780_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1332_ net28 _0170_ _0642_ _0647_ _1332_/VDD _1332_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput5 wbs_adr_i[0] net5 input5/VDD input5/VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_1401_ _0016_ net68 mprj.PS_R1_inst1.LUT_inst1.i3 _1401_/VDD _1401_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1263_ _0576_ _0592_ _0593_ _0594_ _1352_/VDD _1263_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0978_ _0295_ _0322_ _0978_/VDD _0978_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_1246_ _0562_ _0577_ _0103_ _0578_ _1246_/VDD _1246_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0901_ _0244_ _0246_ _0247_ _0901_/VDD _0901_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0694_ net8 _0040_ _0050_ _0694_/VDD _0694_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_0763_ _0112_ _0113_ _0114_ _0115_ _0763_/VDD _0763_/VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_1177_ _0127_ _0385_ _0411_ _0513_ _1177_/VDD _1177_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0832_ _0093_ _0119_ _0130_ _0181_ _0832_/VDD _0832_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1315_ net14 _0637_ _0638_ _1315_/VDD _1315_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1100_ _0367_ _0406_ _0438_ _0439_ _1100_/VDD _1100_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_0746_ _0098_ _0099_ _0746_/VDD _0746_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
Xinput30 wbs_stb_i net30 input30/VDD input30/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_1031_ mprj.PS_Rx_inst7.LUT_inst1.i3 _0373_ _1031_/VDD _1031_/VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_0815_ _0140_ _0162_ _0164_ _0165_ _0815_/VDD _1199_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_0677_ _0032_ _0034_ net35 _0677_/VDD _0677_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1229_ _0546_ _0554_ _0561_ _0562_ _1229_/VDD _1229_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_1014_ _0340_ _0355_ _0356_ _0357_ _1014_/VDD _1014_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0729_ _0078_ _0067_ _0082_ _0083_ _0729_/VDD _0729_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xuser_project_wrapper_208 la_data_out[63] user_project_wrapper_208/VDD user_project_wrapper_208/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0994_ _0336_ _0337_ _0994_/VDD _0994_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1331_ _0646_ _0007_ _1331_/VDD _1331_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1400_ _0015_ net69 mprj.PS_R1_inst1.LUT_inst15.I1 _1400_/VDD _1400_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_1193_ _0190_ _0323_ _0334_ _0528_ _1193_/VDD _1193_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0977_ mprj.PS_Rx_inst7.LUT_inst1.i3 _0295_ _0321_ _1152_/VDD _0977_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xinput6 wbs_adr_i[1] net6 input6/VDD input6/VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_1262_ _0576_ _0592_ _0050_ _0593_ _1262_/VDD _1262_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0831_ _0126_ _0076_ _0138_ _0106_ _0179_ _0180_ _0831_/VDD _0831_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0693_ _0046_ _0048_ _0049_ _0693_/VDD _0693_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1176_ _0491_ _0497_ _0511_ _0512_ _1176_/VDD _1176_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_1314_ _0636_ _0637_ _1314_/VDD _1314_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_0762_ mprj.PS_Rx_inst2.LUT_inst1.i4 mprj.PS_Rx_inst3.LUT_inst1.i3 _0114_ _0762_/VDD
+ _0762_/VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
X_1245_ _0567_ _0576_ _0577_ _1245_/VDD _1245_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_4
X_0900_ _0242_ _0245_ _0246_ _0900_/VDD _0900_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0814_ _0107_ _0076_ _0138_ _0093_ _0163_ _0164_ _0814_/VDD _0814_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1030_ _0070_ _0319_ _0372_ _1030_/VDD _1030_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xinput20 wbs_dat_i[15] net20 input20/VDD input20/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput31 wbs_we_i net31 input31/VDD input31/VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_0745_ _0046_ _0065_ mprj.PS_Rx_inst2.LUT_inst1.i4 _0098_ _0745_/VDD _0745_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1159_ _0494_ _0495_ _0421_ net46 _1159_/VDD _1159_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0676_ net31 net13 net30 _0033_ _0034_ _0676_/VDD _0676_/VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_1228_ _0545_ _0556_ _0560_ _0561_ _1228_/VDD _1228_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_1013_ _0340_ _0355_ _0102_ _0356_ _1013_/VDD _1013_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0728_ _0078_ _0079_ _0081_ _0082_ _0728_/VDD _0728_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xuser_project_wrapper_209 user_irq[0] user_project_wrapper_209/VDD user_project_wrapper_209/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0993_ _0316_ _0335_ _0336_ _0993_/VDD _0993_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1330_ net27 _0147_ _0642_ _0646_ _1330_/VDD _1330_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1261_ _0580_ _0591_ _0592_ _1261_/VDD _1261_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
Xinput7 wbs_adr_i[2] net7 input7/VDD input7/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_0976_ _0319_ _0320_ _0976_/VDD _0976_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1192_ _0510_ _0524_ _0526_ _0527_ _1192_/VDD _1192_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_0830_ _0126_ _0081_ _0099_ _0179_ _0830_/VDD _0830_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0761_ mprj.PS_Rx_inst2.LUT_inst1.i4 mprj.PS_Rx_inst3.LUT_inst1.i3 _0113_ _0761_/VDD
+ _0761_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1244_ _0561_ _0569_ _0575_ _0576_ _1244_/VDD _1244_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_1313_ _0039_ _0635_ _0636_ _1313_/VDD _1313_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_0692_ _0035_ mprj.PS_R1_inst1.LUT_inst1.i1 _0047_ _0048_ _0692_/VDD _0692_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1175_ _0490_ _0499_ _0510_ _0511_ _1175_/VDD _1175_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_0959_ _0070_ _0289_ _0302_ _0303_ _0959_/VDD _0959_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0744_ _0067_ _0073_ _0074_ _0097_ _0744_/VDD _0744_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1158_ _0468_ _0493_ _0103_ _0495_ _1158_/VDD _1158_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0813_ _0106_ _0081_ _0099_ _0163_ _0813_/VDD _0813_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1089_ mprj.PS_R1_inst1.LUT_inst13.I1 _0115_ _0132_ mprj.PS_R1_inst1.LUT_inst12.I1
+ _0427_ _0428_ _1089_/VDD _1089_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xinput10 wbs_adr_i[5] net10 input10/VDD input10/VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput21 wbs_dat_i[1] net21 input21/VDD input21/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_0675_ net6 net5 net8 _0033_ _0675_/VDD _0675_/VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1227_ _0055_ _0543_ _0559_ _0560_ _1227_/VDD _1227_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1012_ _0315_ _0354_ _0355_ _1012_/VDD _1012_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_0727_ _0080_ _0081_ _0727_/VDD _0727_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0992_ _0295_ _0317_ _0335_ _0992_/VDD _0992_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1260_ _0575_ _0582_ _0590_ _0591_ _1260_/VDD _1260_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_1191_ _0240_ _0248_ _0287_ _0217_ _0525_ _0526_ _1191_/VDD _1191_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xinput8 wbs_adr_i[3] net8 input8/VDD input8/VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_0975_ _0316_ _0318_ _0319_ _0975_/VDD _0975_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_1389_ _0004_ net70 mprj.PS_R1_inst1.LUT_inst4.I1 _1389_/VDD _1389_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0760_ _0104_ _0112_ _0760_/VDD _0760_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_0691_ mprj.PS_R1_inst1.LUT_inst1.i3 _0047_ _0691_/VDD _0691_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_1312_ net4 net2 _0034_ _0635_ _1312_/VDD _1312_/VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1174_ _0487_ _0502_ _0509_ _0510_ _1174_/VDD _1174_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_0889_ _0225_ _0234_ _0103_ _0236_ _0889_/VDD _0889_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0958_ _0070_ _0248_ _0287_ _0301_ _0302_ _0958_/VDD _0958_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
Xuser_project_wrapper_190 la_data_out[45] user_project_wrapper_190/VDD user_project_wrapper_190/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1243_ _0560_ _0572_ _0574_ _0575_ _1243_/VDD _1243_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1226_ _0449_ _0220_ _0557_ _0558_ _0559_ _1226_/VDD _1226_/VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_0812_ _0070_ _0130_ _0160_ _0161_ _0162_ _0812_/VDD _0812_/VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_0674_ net10 net9 net12 net11 _0032_ _0674_/VDD _0674_/VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_0743_ _0065_ _0067_ _0059_ _0096_ _0743_/VDD _0743_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xinput11 wbs_adr_i[6] net11 input11/VDD input11/VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput22 wbs_dat_i[2] net22 input22/VDD input22/VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_1157_ _0468_ _0493_ _0494_ _1157_/VDD _1157_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
X_1088_ mprj.PS_R1_inst1.LUT_inst13.I1 _0119_ _0130_ _0427_ _1088_/VDD _1088_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1011_ _0314_ _0342_ _0353_ _0354_ _1011_/VDD _1011_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1209_ _0155_ _0540_ _0542_ _0543_ _1209_/VDD _1209_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0726_ mprj.PS_R1_inst1.LUT_inst1.i4 mprj.PS_Rx_inst2.LUT_inst1.i3 _0080_ _0726_/VDD
+ _0726_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_0709_ _0060_ _0064_ _0709_/VDD _0709_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0991_ _0333_ _0334_ _0991_/VDD _0991_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1190_ _0239_ _0249_ _0289_ _0525_ _1190_/VDD _1190_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xinput9 wbs_adr_i[4] net9 input9/VDD input9/VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_0974_ _0295_ _0317_ _0318_ _0974_/VDD _0974_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1388_ _0003_ net68 mprj.PS_R1_inst1.LUT_inst3.I1 _1388_/VDD _1388_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0690_ mprj.PS_R1_inst1.LUT_inst1.i4 _0046_ _0690_/VDD _1132_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0888_ _0225_ _0234_ _0235_ _0888_/VDD _0888_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1173_ _0506_ _0508_ _0509_ _1173_/VDD _1173_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1311_ net1 net34 _1311_/VDD _1311_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1242_ _0330_ _0248_ _0287_ _0298_ _0573_ _0574_ _1242_/VDD _1242_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0957_ _0300_ _0301_ _0957_/VDD _0957_/VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xuser_project_wrapper_180 la_data_out[35] user_project_wrapper_180/VDD user_project_wrapper_180/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_191 la_data_out[46] user_project_wrapper_191/VDD user_project_wrapper_191/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0811_ mprj.PS_R1_inst1.LUT_inst2.I1 _0117_ _0132_ _0161_ _0811_/VDD _0811_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0742_ net8 _0094_ _0040_ _0095_ _0742_/VDD _0742_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xinput12 wbs_adr_i[7] net12 input12/VDD input12/VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput23 wbs_dat_i[3] net23 input8/VDD input23/VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_1156_ _0475_ _0492_ _0493_ _1156_/VDD _1156_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_1225_ _0330_ _0206_ _0222_ _0558_ _1225_/VDD _1225_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1087_ _0046_ _0425_ _0426_ _1087_/VDD _1087_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_1010_ _0313_ _0344_ _0352_ _0353_ _1010_/VDD _1010_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_1208_ _0112_ _0449_ _0541_ _0330_ _0154_ _0542_ _1208_/VDD _1208_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1139_ _0147_ _0323_ _0334_ _0476_ _1139_/VDD _1139_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0725_ mprj.PS_R1_inst1.LUT_inst1.i4 _0065_ _0079_ _0725_/VDD _0725_/VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
X_0708_ _0062_ _0063_ _0708_/VDD _0708_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0990_ _0237_ mprj.PS_Rx_inst7.LUT_inst1.i3 _0295_ _0333_ _0990_/VDD _0990_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1387_ _0002_ net70 mprj.PS_R1_inst1.LUT_inst2.I1 _1387_/VDD _1387_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0973_ _0237_ mprj.PS_Rx_inst7.LUT_inst1.i3 _0317_ _0973_/VDD _0973_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1310_ _0051_ _0055_ _0421_ net60 _1310_/VDD _1310_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0956_ mprj.PS_Rx_inst6.LUT_inst1.i3 _0237_ mprj.PS_R1_inst1.LUT_inst2.I1 _0300_
+ _0956_/VDD _0956_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1172_ _0269_ _0204_ _0221_ _0239_ _0507_ _0508_ _1172_/VDD _1172_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1241_ _0330_ _0249_ _0289_ _0573_ _1241_/VDD _1241_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0887_ _0200_ _0233_ _0234_ _0887_/VDD _0887_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
Xuser_project_wrapper_170 la_data_out[25] user_project_wrapper_170/VDD user_project_wrapper_170/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_181 la_data_out[36] user_project_wrapper_181/VDD user_project_wrapper_181/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_192 la_data_out[47] user_project_wrapper_192/VDD user_project_wrapper_192/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0810_ _0070_ _0116_ _0160_ _0810_/VDD _0810_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xinput24 wbs_dat_i[4] net24 input24/VDD input24/VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput13 wbs_cyc_i net13 input13/VDD input13/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_0741_ _0093_ _0094_ _0741_/VDD _1384_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1086_ mprj.PS_R1_inst1.LUT_inst15.I1 _0075_ _0138_ mprj.PS_R1_inst1.LUT_inst14.I1
+ _0424_ _0425_ _1086_/VDD _1086_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1155_ _0467_ _0477_ _0491_ _0492_ _1155_/VDD _1155_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1224_ _0449_ _0205_ _0557_ _1224_/VDD _1224_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_0939_ _0283_ _0284_ _0939_/VDD _0939_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_0724_ mprj.PS_R1_inst1.LUT_inst1.i0 _0078_ _0724_/VDD _0724_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1207_ _0112_ mprj.PS_Rx_inst4.LUT_inst1.i3 _0541_ _1207_/VDD _1207_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1069_ _0371_ _0394_ _0408_ _0409_ _1069_/VDD _1069_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1138_ _0107_ _0382_ _0443_ _0094_ _0474_ _0475_ _1138_/VDD _1138_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0707_ mprj.PS_R1_inst1.LUT_inst2.I1 _0062_ _0707_/VDD _0707_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1386_ _0001_ net70 mprj.PS_R1_inst1.LUT_inst1.i1 _1386_/VDD _1386_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0972_ _0237_ mprj.PS_Rx_inst7.LUT_inst1.i3 _0316_ _0972_/VDD _0972_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1240_ _0390_ _0203_ _0570_ _0571_ _0572_ _1240_/VDD _1240_/VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_1171_ _0269_ _0209_ _0219_ _0507_ _1171_/VDD _1171_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0955_ _0058_ _0298_ _0060_ _0299_ _0955_/VDD _0955_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1369_ net29 _0657_ _0667_ _1369_/VDD _1369_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xuser_project_wrapper_160 la_data_out[15] user_project_wrapper_160/VDD user_project_wrapper_160/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_171 la_data_out[26] user_project_wrapper_171/VDD user_project_wrapper_171/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_182 la_data_out[37] user_project_wrapper_182/VDD user_project_wrapper_182/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_193 la_data_out[48] user_project_wrapper_193/VDD user_project_wrapper_193/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0886_ _0199_ _0230_ _0232_ _0233_ _0886_/VDD _0886_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_0740_ mprj.PS_R1_inst1.LUT_inst4.I1 _0093_ _0740_/VDD _0740_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xinput25 wbs_dat_i[5] net25 input25/VDD input25/VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput14 wbs_dat_i[0] net14 input14/VDD input14/VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_0869_ mprj.PS_R1_inst1.LUT_inst10.I1 _0216_ _0869_/VDD _0869_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1085_ mprj.PS_R1_inst1.LUT_inst15.I1 _0080_ _0098_ _0424_ _1085_/VDD _1085_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1223_ _0298_ _0248_ _0287_ _0270_ _0555_ _0556_ _1223_/VDD _1223_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0938_ mprj.PS_Rx_inst6.LUT_inst1.i3 _0237_ mprj.PS_R1_inst1.LUT_inst1.i1 _0283_
+ _0938_/VDD _0938_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1154_ _0463_ _0479_ _0490_ _0491_ _1154_/VDD _1154_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_0723_ mprj.PS_R1_inst1.LUT_inst1.i1 _0076_ _0077_ _0723_/VDD _0723_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1206_ _0144_ _0390_ _0540_ _1206_/VDD _1206_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1137_ _0107_ _0385_ _0411_ _0474_ _1137_/VDD _1137_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1068_ _0370_ _0396_ _0407_ _0408_ _1068_/VDD _1068_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_0706_ _0049_ _0051_ _0055_ _0056_ _0061_ net47 _0706_/VDD _0706_/VSS gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_0971_ _0282_ _0303_ _0314_ _0315_ _0971_/VDD _0971_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_1385_ _0000_ net71 mprj.PS_R1_inst1.LUT_inst1.i0 _1385_/VDD _1385_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_1170_ _0503_ _0504_ _0505_ _0506_ _1170_/VDD _1170_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0885_ _0093_ _0157_ _0175_ mprj.PS_R1_inst1.LUT_inst3.I1 _0231_ _0232_ _0885_/VDD
+ _0885_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1299_ _0586_ _0382_ _0626_ _1299_/VDD _1299_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0954_ _0297_ _0298_ _0954_/VDD _0954_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
Xuser_project_wrapper_161 la_data_out[16] user_project_wrapper_161/VDD user_project_wrapper_161/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_150 la_data_out[5] user_project_wrapper_150/VDD user_project_wrapper_150/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_172 la_data_out[27] user_project_wrapper_172/VDD user_project_wrapper_172/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_183 la_data_out[38] user_project_wrapper_183/VDD user_project_wrapper_183/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_194 la_data_out[49] user_project_wrapper_194/VDD user_project_wrapper_194/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1368_ _0666_ _0024_ _1368_/VDD _1368_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1222_ _0297_ _0249_ _0289_ _0555_ _1222_/VDD _1222_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1084_ _0107_ _0320_ _0337_ _0094_ _0422_ _0423_ _1084_/VDD _1084_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1153_ _0460_ _0487_ _0489_ _0490_ _1153_/VDD _1153_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_2
Xinput15 wbs_dat_i[10] net15 input15/VDD input15/VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput26 wbs_dat_i[6] net26 input26/VDD input26/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0868_ mprj.PS_Rx_inst6.LUT_inst1.i3 _0068_ _0215_ _0868_/VDD _0868_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0799_ mprj.PS_Rx_inst4.LUT_inst1.i3 _0144_ _0149_ _0799_/VDD _0799_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_0937_ _0261_ _0273_ _0281_ _0282_ _0937_/VDD _0937_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_0722_ _0075_ _0076_ _0722_/VDD _0722_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1136_ _0472_ _0473_ _0421_ net45 _1136_/VDD _1136_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1067_ _0367_ _0404_ _0406_ _0407_ _1067_/VDD _1067_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1205_ _0330_ _0204_ _0221_ _0297_ _0538_ _0539_ _1205_/VDD _1205_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0705_ _0058_ _0059_ _0060_ _0061_ _0705_/VDD _0705_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1119_ _0454_ _0456_ _0457_ _1119_/VDD _1119_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_0970_ _0281_ _0305_ _0313_ _0314_ _0970_/VDD _0970_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_1384_ mprj.PS_Rx_inst8.carry_inst.O net68 net33 _1384_/VDD _1384_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1367_ net28 mprj.PS_Rx_inst5.LUT_inst1.i3 _0655_ _0666_ _1367_/VDD _1367_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0953_ mprj.PS_R1_inst1.LUT_inst13.I1 _0297_ _0953_/VDD _0953_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0884_ _0093_ _0152_ _0173_ _0231_ _0884_/VDD _0884_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xuser_project_wrapper_162 la_data_out[17] user_project_wrapper_162/VDD user_project_wrapper_162/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_151 la_data_out[6] user_project_wrapper_151/VDD user_project_wrapper_151/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_173 la_data_out[28] user_project_wrapper_173/VDD user_project_wrapper_173/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_184 la_data_out[39] user_project_wrapper_184/VDD user_project_wrapper_184/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_195 la_data_out[50] user_project_wrapper_195/VDD user_project_wrapper_195/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_140 io_out[33] user_project_wrapper_140/VDD user_project_wrapper_140/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1298_ _0331_ _0383_ _0443_ _0625_ _1298_/VDD _1298_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1152_ _0239_ _0205_ _0222_ _0216_ _0488_ _0489_ _1152_/VDD _1152_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1083_ _0107_ _0323_ _0334_ _0422_ _1083_/VDD _1083_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1221_ _0240_ _0319_ _0336_ _0217_ _0553_ _0554_ _1221_/VDD _1221_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xinput16 wbs_dat_i[11] net16 input16/VDD input16/VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput27 wbs_dat_i[7] net27 input27/VDD input27/VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_0936_ _0260_ _0275_ _0280_ _0281_ _0936_/VDD _0936_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_0867_ _0188_ _0191_ _0214_ net67 _0867_/VDD _0867_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0798_ _0058_ _0147_ _0064_ _0148_ _0798_/VDD _0798_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1066_ _0169_ _0205_ _0222_ _0146_ _0405_ _0406_ _1066_/VDD _1066_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1204_ _0330_ _0208_ _0219_ _0538_ _1204_/VDD _1204_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0721_ mprj.PS_Rx_inst2.LUT_inst1.i4 _0073_ _0074_ _0075_ _0721_/VDD _0721_/VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1135_ _0468_ _0471_ _0103_ _0473_ _1135_/VDD _1135_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0919_ _0233_ _0261_ _0264_ _0265_ _0919_/VDD _0919_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_0704_ _0036_ _0038_ _0039_ _0060_ _0704_/VDD _0704_/VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_1118_ mprj.PS_R1_inst1.LUT_inst14.I1 _0116_ _0132_ _0297_ _0455_ _0456_ _1118_/VDD
+ _1118_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1049_ mprj.PS_R1_inst1.LUT_inst15.I1 _0390_ _1049_/VDD _1049_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_1383_ mprj.PS_R1_inst1.LUT_inst1.i0 net71 net32 _1383_/VDD _1383_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xuser_project_wrapper_130 io_out[23] user_project_wrapper_130/VDD user_project_wrapper_130/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0883_ _0196_ _0227_ _0229_ _0230_ _0883_/VDD _0883_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_0952_ _0295_ _0068_ _0296_ _0952_/VDD _0952_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xuser_project_wrapper_163 la_data_out[18] user_project_wrapper_163/VDD user_project_wrapper_163/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_152 la_data_out[7] user_project_wrapper_152/VDD user_project_wrapper_152/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_174 la_data_out[29] user_project_wrapper_174/VDD user_project_wrapper_174/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_141 io_out[34] user_project_wrapper_141/VDD user_project_wrapper_141/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1366_ _0154_ _0656_ _0665_ _0023_ _1366_/VDD _1366_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xuser_project_wrapper_185 la_data_out[40] user_project_wrapper_185/VDD user_project_wrapper_185/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_196 la_data_out[51] user_project_wrapper_196/VDD user_project_wrapper_196/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1297_ _0421_ _0624_ net56 _1297_/VDD _1297_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1151_ _0239_ _0209_ _0220_ _0488_ _1151_/VDD _1151_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1220_ _0240_ _0323_ _0333_ _0553_ _1220_/VDD _1220_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xinput17 wbs_dat_i[12] net17 input17/VDD input17/VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput28 wbs_dat_i[8] net28 input28/VDD input28/VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_0935_ _0259_ _0277_ _0279_ _0280_ _0935_/VDD _0935_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_0866_ _0200_ _0212_ _0213_ _0214_ _0866_/VDD _0866_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1349_ _0655_ _0656_ _1349_/VDD _1349_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1082_ _0418_ _0419_ _0421_ net43 _1082_/VDD _1082_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0797_ _0146_ _0147_ _0797_/VDD _0797_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1203_ _0270_ _0248_ _0287_ _0240_ _0536_ _0537_ _1203_/VDD _1203_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1065_ _0169_ _0209_ _0220_ _0405_ _1065_/VDD _1065_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0720_ _0046_ _0065_ _0074_ _0720_/VDD _0720_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
X_1134_ _0468_ _0471_ _0472_ _1134_/VDD _1134_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
X_0918_ _0071_ _0220_ _0262_ _0263_ _0264_ _0918_/VDD _0918_/VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_0849_ _0106_ _0119_ _0130_ _0197_ _0849_/VDD _0849_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0703_ mprj.PS_R1_inst1.LUT_inst1.i1 _0059_ _0703_/VDD _0703_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1117_ mprj.PS_R1_inst1.LUT_inst14.I1 _0119_ _0130_ _0455_ _1117_/VDD _1117_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1048_ _0103_ mprj.PS_Rx_inst8.carry_inst.O _0389_ _1048_/VDD _1048_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1382_ _0673_ _0031_ _1382_/VDD _1382_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0951_ mprj.PS_Rx_inst7.LUT_inst1.i4 _0295_ _0951_/VDD _0951_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0882_ _0169_ _0075_ _0137_ mprj.PS_R1_inst1.LUT_inst7.I1 _0228_ _0229_ _0882_/VDD
+ _0882_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xuser_project_wrapper_131 io_out[24] user_project_wrapper_131/VDD user_project_wrapper_131/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_120 io_out[13] user_project_wrapper_120/VDD user_project_wrapper_120/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_153 la_data_out[8] user_project_wrapper_153/VDD user_project_wrapper_153/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_164 la_data_out[19] user_project_wrapper_164/VDD user_project_wrapper_164/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_175 la_data_out[30] user_project_wrapper_175/VDD user_project_wrapper_175/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_186 la_data_out[41] user_project_wrapper_186/VDD user_project_wrapper_186/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_197 la_data_out[52] user_project_wrapper_197/VDD user_project_wrapper_197/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_142 io_out[35] user_project_wrapper_142/VDD user_project_wrapper_142/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1365_ net27 _0657_ _0665_ _1365_/VDD _1365_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1296_ _0612_ _0622_ _0623_ _0624_ _1296_/VDD _1296_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xinput18 wbs_dat_i[13] net18 input18/VDD input18/VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput29 wbs_dat_i[9] net29 input29/VDD input29/VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_0934_ mprj.PS_R1_inst1.LUT_inst10.I1 _0075_ _0138_ mprj.PS_R1_inst1.LUT_inst10.I0
+ _0278_ _0279_ _0934_/VDD _0934_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0865_ _0200_ _0212_ _0050_ _0213_ _0865_/VDD _0865_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0796_ mprj.PS_R1_inst1.LUT_inst7.I1 _0146_ _0796_/VDD _0796_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1081_ _0420_ _0421_ _1081_/VDD _1081_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1150_ _0457_ _0482_ _0486_ _0487_ _1150_/VDD _1150_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1348_ _0042_ _0635_ _0655_ _1348_/VDD _1348_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1279_ _0298_ _0381_ _0413_ _0270_ _0607_ _0608_ _1279_/VDD _1279_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1133_ _0441_ _0470_ _0471_ _1133_/VDD _1133_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1202_ _0269_ _0249_ _0289_ _0536_ _1202_/VDD _1202_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1064_ _0366_ _0398_ _0403_ _0404_ _1064_/VDD _1064_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_0779_ _0129_ _0130_ _0779_/VDD _0779_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_0848_ _0146_ _0076_ _0138_ _0126_ _0195_ _0196_ _0848_/VDD _0848_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0917_ _0062_ _0206_ _0222_ _0263_ _0917_/VDD _0917_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0702_ _0057_ _0058_ _0702_/VDD _0702_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1047_ _0388_ mprj.PS_Rx_inst8.carry_inst.O _1047_/VDD _1047_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1116_ _0073_ _0450_ _0452_ _0453_ _0454_ _1116_/VDD _1116_/VSS gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_1381_ net20 mprj.PS_Rx_inst8.LUT_inst1.i4 _0655_ _0673_ _1381_/VDD _1381_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xuser_project_wrapper_121 io_out[14] user_project_wrapper_121/VDD user_project_wrapper_121/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_132 io_out[25] user_project_wrapper_132/VDD user_project_wrapper_132/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0950_ _0268_ _0271_ _0294_ net39 _0950_/VDD _0950_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1364_ _0664_ _0022_ _1364_/VDD _1364_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0881_ mprj.PS_R1_inst1.LUT_inst8.I1 _0080_ _0098_ _0228_ _0881_/VDD _0881_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xuser_project_wrapper_154 la_data_out[9] user_project_wrapper_154/VDD user_project_wrapper_154/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_165 la_data_out[20] user_project_wrapper_165/VDD user_project_wrapper_165/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_176 la_data_out[31] user_project_wrapper_176/VDD user_project_wrapper_176/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_187 la_data_out[42] user_project_wrapper_187/VDD user_project_wrapper_187/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_198 la_data_out[53] user_project_wrapper_198/VDD user_project_wrapper_198/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_143 io_out[36] user_project_wrapper_143/VDD user_project_wrapper_143/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1295_ _0612_ _0622_ _0050_ _0623_ _1295_/VDD _1295_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xuser_project_wrapper_110 io_out[3] user_project_wrapper_110/VDD user_project_wrapper_110/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput19 wbs_dat_i[14] net19 input19/VDD input19/VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_0864_ _0201_ _0211_ _0212_ _0864_/VDD _0864_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1080_ _0060_ _0043_ _0420_ _1080_/VDD _1080_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_0933_ mprj.PS_R1_inst1.LUT_inst10.I1 _0081_ _0099_ _0278_ _0933_/VDD _0933_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0795_ _0144_ _0068_ _0145_ _0795_/VDD _0795_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1278_ _0298_ _0385_ _0410_ _0607_ _1278_/VDD _1278_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1416_ _0031_ net71 mprj.PS_Rx_inst8.LUT_inst1.i4 _1416_/VDD _1416_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_1347_ _0390_ _0637_ _0654_ _0015_ _1347_/VDD _1347_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1201_ _0217_ _0319_ _0336_ _0190_ _0534_ _0535_ _1201_/VDD _1201_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1132_ _0094_ _0382_ _0443_ _0071_ _0469_ _0470_ _1132_/VDD _1132_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0916_ _0071_ _0205_ _0262_ _0916_/VDD _0916_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0778_ mprj.PS_Rx_inst2.LUT_inst1.i4 mprj.PS_Rx_inst3.LUT_inst1.i3 _0104_ _0129_
+ _0778_/VDD _0778_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0847_ _0146_ _0081_ _0099_ _0195_ _0847_/VDD _0847_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1063_ _0365_ _0400_ _0402_ _0403_ _1063_/VDD _1063_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_1115_ _0046_ _0390_ _0067_ _0453_ _1115_/VDD _1115_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1046_ mprj.PS_Rx_inst8.LUT_inst1.i4 _0377_ _0387_ _0388_ _1046_/VDD _1046_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_0701_ net8 _0057_ _0701_/VDD _0701_/VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_1029_ _0353_ _0359_ _0370_ _0371_ _1029_/VDD _1029_/VSS gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_1380_ _0672_ _0030_ _1380_/VDD _1380_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xuser_project_wrapper_122 io_out[15] user_project_wrapper_122/VDD user_project_wrapper_122/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1294_ _0617_ _0621_ _0622_ _1294_/VDD _1294_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
Xuser_project_wrapper_133 io_out[26] user_project_wrapper_133/VDD user_project_wrapper_133/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0880_ _0126_ _0116_ _0132_ mprj.PS_R1_inst1.LUT_inst5.I1 _0226_ _0227_ _0880_/VDD
+ _0880_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xuser_project_wrapper_100 io_oeb[28] user_project_wrapper_100/VDD user_project_wrapper_100/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_111 io_out[4] user_project_wrapper_111/VDD user_project_wrapper_111/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_155 la_data_out[10] user_project_wrapper_155/VDD user_project_wrapper_155/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_166 la_data_out[21] user_project_wrapper_166/VDD user_project_wrapper_166/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_177 la_data_out[32] user_project_wrapper_177/VDD user_project_wrapper_177/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_188 la_data_out[43] user_project_wrapper_188/VDD user_project_wrapper_188/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_199 la_data_out[54] user_project_wrapper_199/VDD user_project_wrapper_199/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_144 io_out[37] user_project_wrapper_144/VDD user_project_wrapper_144/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1363_ net26 mprj.PS_Rx_inst4.LUT_inst1.i3 _0655_ _0664_ _1363_/VDD _1363_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0932_ mprj.PS_R1_inst1.LUT_inst8.I1 _0115_ _0131_ mprj.PS_R1_inst1.LUT_inst7.I1
+ _0276_ _0277_ _0932_/VDD _0932_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1277_ _0605_ _0606_ _0421_ net54 _1277_/VDD _1277_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0863_ _0059_ _0205_ _0210_ _0211_ _0863_/VDD _0863_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0794_ mprj.PS_Rx_inst4.LUT_inst1.i4 _0144_ _1010_/VDD _0794_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1415_ _0030_ net68 mprj.PS_Rx_inst8.LUT_inst1.i3 _1415_/VDD _1415_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_1346_ net20 _0637_ _0654_ _1346_/VDD _1346_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0915_ _0230_ _0255_ _0260_ _0261_ _0915_/VDD _0915_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1062_ mprj.PS_R1_inst1.LUT_inst14.I1 _0075_ _0138_ mprj.PS_R1_inst1.LUT_inst13.I1
+ _0401_ _0402_ _1062_/VDD _1062_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1131_ _0094_ _0385_ _0411_ _0469_ _1131_/VDD _1131_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0777_ _0058_ _0127_ _0064_ _0128_ _0777_/VDD _0777_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1200_ _0217_ _0316_ _0333_ _0534_ _1200_/VDD _1200_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0846_ _0071_ _0173_ _0192_ _0193_ _0194_ _0846_/VDD _0846_/VSS gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1329_ _0645_ _0006_ _1329_/VDD _1329_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0700_ _0046_ _0043_ _0056_ _0700_/VDD _0700_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1114_ _0052_ _0065_ _0451_ _0452_ _1114_/VDD _1114_/VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1045_ mprj.PS_R1_inst1.LUT_inst1.i1 _0382_ _0384_ _0386_ _0387_ _1045_/VDD _1045_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_0829_ _0063_ _0173_ _0176_ _0177_ _0178_ _0829_/VDD _0829_/VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1028_ _0352_ _0367_ _0369_ _0370_ _1028_/VDD _1028_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
Xuser_project_wrapper_123 io_out[16] user_project_wrapper_123/VDD user_project_wrapper_123/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1293_ _0603_ _0620_ _0621_ _1293_/VDD _1293_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xuser_project_wrapper_134 io_out[27] user_project_wrapper_134/VDD user_project_wrapper_134/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_101 io_oeb[29] user_project_wrapper_101/VDD user_project_wrapper_101/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_112 io_out[5] user_project_wrapper_112/VDD user_project_wrapper_112/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_156 la_data_out[11] user_project_wrapper_156/VDD user_project_wrapper_156/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_145 la_data_out[0] user_project_wrapper_145/VDD user_project_wrapper_145/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_167 la_data_out[22] user_project_wrapper_167/VDD user_project_wrapper_167/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_178 la_data_out[33] user_project_wrapper_178/VDD user_project_wrapper_178/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_189 la_data_out[44] user_project_wrapper_189/VDD user_project_wrapper_189/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1362_ _0112_ _0656_ _0663_ _0021_ _1362_/VDD _1362_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0793_ _0125_ _0128_ _0142_ _0143_ net64 _0793_/VDD _0793_/VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_0862_ _0078_ _0144_ _0206_ _0207_ _0209_ _0210_ _0862_/VDD _0862_/VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_1345_ _0451_ _0637_ _0653_ _0014_ _1345_/VDD _1345_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0931_ mprj.PS_R1_inst1.LUT_inst8.I1 _0113_ _0129_ _0276_ _0931_/VDD _0931_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1414_ _0029_ net68 mprj.PS_Rx_inst7.LUT_inst1.i4 _1414_/VDD _1414_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1276_ _0591_ _0604_ _0103_ _0606_ _1276_/VDD _1276_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1061_ mprj.PS_R1_inst1.LUT_inst14.I1 _0081_ _0098_ _0401_ _1061_/VDD _1061_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1130_ _0440_ _0448_ _0467_ _0468_ _1130_/VDD _1130_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_0845_ mprj.PS_R1_inst1.LUT_inst2.I1 _0149_ _0175_ _0193_ _0845_/VDD _0845_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0914_ _0229_ _0257_ _0259_ _0260_ _0914_/VDD _0914_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_1328_ net26 _0127_ _0642_ _0645_ _1328_/VDD _1328_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1259_ _0086_ _0572_ _0589_ _0590_ _1259_/VDD _1259_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_0776_ _0126_ _0127_ _0776_/VDD _0776_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0828_ _0062_ _0157_ _0177_ _0828_/VDD _0828_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1113_ mprj.PS_R1_inst1.LUT_inst14.I1 _0451_ _1113_/VDD _1113_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_1044_ _0078_ _0383_ _0385_ _0386_ _1044_/VDD _1044_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0759_ _0071_ _0076_ _0110_ _0111_ _0759_/VDD _0759_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1027_ _0146_ _0205_ _0222_ _0126_ _0368_ _0369_ _1027_/VDD _1027_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xuser_project_wrapper_124 io_out[17] user_project_wrapper_124/VDD user_project_wrapper_124/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_135 io_out[28] user_project_wrapper_135/VDD user_project_wrapper_135/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_102 io_oeb[30] user_project_wrapper_102/VDD user_project_wrapper_102/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_113 io_out[6] user_project_wrapper_113/VDD user_project_wrapper_113/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_157 la_data_out[12] user_project_wrapper_157/VDD user_project_wrapper_157/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_146 la_data_out[1] user_project_wrapper_146/VDD user_project_wrapper_146/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_168 la_data_out[23] user_project_wrapper_168/VDD user_project_wrapper_168/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_179 la_data_out[34] user_project_wrapper_179/VDD user_project_wrapper_179/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1361_ net25 _0657_ _0663_ _1361_/VDD _1361_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1292_ _0586_ _0318_ _0618_ _0619_ _0620_ _1292_/VDD _1292_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_1275_ _0591_ _0604_ _0605_ _1275_/VDD _1275_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
X_0792_ _0135_ _0141_ _0103_ _0143_ _0792_/VDD _0792_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1413_ _0028_ net69 mprj.PS_Rx_inst7.LUT_inst1.i3 _1413_/VDD _1413_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_1344_ net19 _0637_ _0653_ _1344_/VDD _1344_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_0930_ mprj.PS_R1_inst1.LUT_inst6.I1 _0156_ _0174_ mprj.PS_R1_inst1.LUT_inst5.I1
+ _0274_ _0275_ _0930_/VDD _0930_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0861_ _0208_ _0209_ _0861_/VDD _0861_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1060_ _0269_ _0116_ _0132_ mprj.PS_R1_inst1.LUT_inst11.I1 _0399_ _0400_ _1060_/VDD
+ _1060_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0775_ mprj.PS_R1_inst1.LUT_inst6.I1 _0126_ _0775_/VDD _0775_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0844_ _0070_ _0157_ _0192_ _0844_/VDD _0844_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1189_ _0502_ _0519_ _0523_ _0524_ _1189_/VDD _1189_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1258_ _0584_ _0588_ _0589_ _1258_/VDD _1258_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1327_ _0644_ _0005_ _1327_/VDD _1327_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0913_ mprj.PS_R1_inst1.LUT_inst10.I0 _0075_ _0137_ mprj.PS_R1_inst1.LUT_inst8.I1
+ _0258_ _0259_ _0913_/VDD _0913_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1043_ _0378_ _0385_ _1043_/VDD _1043_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1112_ _0136_ _0449_ _0450_ _1112_/VDD _1112_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0758_ _0071_ _0099_ _0109_ _0097_ _0110_ _0758_/VDD _0758_/VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_0827_ _0059_ _0149_ _0175_ _0176_ _0827_/VDD _0827_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0689_ _0035_ _0040_ _0044_ _0045_ net36 _0689_/VDD _0689_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1026_ _0146_ _0209_ _0220_ _0368_ _1026_/VDD _1026_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1009_ _0312_ _0346_ _0351_ _0352_ _1009_/VDD _1009_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
Xuser_project_wrapper_125 io_out[18] user_project_wrapper_125/VDD user_project_wrapper_125/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1291_ _0242_ _0586_ _0322_ _0619_ _1291_/VDD _1291_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xuser_project_wrapper_136 io_out[29] user_project_wrapper_136/VDD user_project_wrapper_136/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_114 io_out[7] user_project_wrapper_114/VDD user_project_wrapper_114/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_103 io_oeb[31] user_project_wrapper_103/VDD user_project_wrapper_103/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_158 la_data_out[13] user_project_wrapper_158/VDD user_project_wrapper_158/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_147 la_data_out[2] user_project_wrapper_147/VDD user_project_wrapper_147/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_169 la_data_out[24] user_project_wrapper_169/VDD user_project_wrapper_169/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1360_ _0662_ _0020_ _1360_/VDD _1360_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0860_ _0144_ mprj.PS_Rx_inst5.LUT_inst1.i3 _0208_ _0860_/VDD _0860_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1343_ _0652_ _0013_ _1343_/VDD _1343_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1412_ _0027_ net71 mprj.PS_Rx_inst6.LUT_inst1.i4 _1412_/VDD _1412_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_0791_ _0135_ _0141_ _0142_ _0791_/VDD _0791_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
X_0989_ net8 _0331_ _0040_ _0332_ _0989_/VDD _0989_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1274_ _0597_ _0599_ _0603_ _0604_ _1274_/VDD _1274_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_1188_ _0055_ _0522_ _0523_ _1188_/VDD _1188_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_0774_ mprj.PS_Rx_inst4.LUT_inst1.i3 _0068_ _0125_ _0774_/VDD _0774_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1257_ _0287_ _0585_ _0587_ _0588_ _1257_/VDD _1257_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0912_ mprj.PS_R1_inst1.LUT_inst10.I0 _0080_ _0098_ _0258_ _0912_/VDD _0912_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0843_ _0058_ _0190_ _0064_ _0191_ _0843_/VDD _0843_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1326_ net25 _0107_ _0642_ _0644_ _1326_/VDD _1326_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1042_ mprj.PS_R1_inst1.LUT_inst1.i0 _0322_ _0383_ _0384_ _1042_/VDD _1042_/VSS gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1111_ mprj.PS_R1_inst1.LUT_inst15.I1 _0449_ _1111_/VDD _1111_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0688_ _0036_ _0039_ mprj.PS_R1_inst1.LUT_inst1.i3 _0045_ _0688_/VDD _0688_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0826_ _0174_ _0175_ _0826_/VDD _0826_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_0757_ _0065_ _0067_ _0062_ _0109_ _0757_/VDD _0757_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1309_ _0421_ _0634_ net59 _1309_/VDD _1309_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0809_ _0144_ _0153_ _0158_ _0159_ _0809_/VDD _0809_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1025_ _0351_ _0361_ _0366_ _0367_ _1025_/VDD _1025_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_1008_ _0311_ _0348_ _0350_ _0351_ _1008_/VDD _1008_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_2
Xuser_project_wrapper_126 io_out[19] user_project_wrapper_126/VDD user_project_wrapper_126/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1290_ _0237_ _0373_ _0331_ _0618_ _1290_/VDD _1290_/VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xuser_project_wrapper_115 io_out[8] user_project_wrapper_115/VDD user_project_wrapper_115/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_137 io_out[30] user_project_wrapper_137/VDD user_project_wrapper_137/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_104 io_oeb[32] user_project_wrapper_104/VDD user_project_wrapper_104/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_159 la_data_out[14] user_project_wrapper_159/VDD user_project_wrapper_159/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_148 la_data_out[3] user_project_wrapper_148/VDD user_project_wrapper_148/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xoutput60 net60 wbs_dat_o[31] output60/VDD output60/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_0790_ _0111_ _0140_ _0141_ _0790_/VDD _0790_/VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1273_ _0601_ _0602_ _0583_ _0603_ _1273_/VDD _1273_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1411_ _0026_ net70 mprj.PS_Rx_inst6.LUT_inst1.i3 _1411_/VDD _1411_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_1342_ net18 _0298_ _0642_ _0652_ _1342_/VDD _1342_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0988_ _0330_ _0331_ _0988_/VDD _0988_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_0911_ mprj.PS_R1_inst1.LUT_inst7.I1 _0115_ _0131_ mprj.PS_R1_inst1.LUT_inst6.I1
+ _0256_ _0257_ _0911_/VDD _0911_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0773_ _0105_ _0108_ _0124_ net63 _0773_/VDD _0773_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1256_ _0586_ _0289_ _0587_ _1256_/VDD _1256_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1325_ _0643_ _0004_ _1325_/VDD _1325_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0842_ _0189_ _0190_ _0842_/VDD _0842_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1187_ _0449_ _0173_ _0520_ _0521_ _0522_ _1187_/VDD _1187_/VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1110_ _0127_ _0320_ _0337_ _0107_ _0447_ _0448_ _1110_/VDD _1110_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1041_ mprj.PS_Rx_inst8.LUT_inst1.i3 mprj.PS_Rx_inst8.LUT_inst1.i4 _0383_ _1041_/VDD
+ _1041_/VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_0756_ _0058_ _0107_ _0064_ _0108_ _0756_/VDD _0756_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0825_ _0154_ _0155_ _0151_ _0174_ _1055_/VDD _0825_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_0687_ _0043_ _0044_ _0687_/VDD _0687_/VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_1308_ _0633_ _0634_ _1308_/VDD _1308_/VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1239_ _0144_ _0390_ _0187_ _0571_ _1239_/VDD _1239_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0808_ _0059_ _0157_ _0153_ _0144_ _0158_ _0808_/VDD _0808_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_1024_ _0350_ _0363_ _0365_ _0366_ _1024_/VDD _1024_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_0739_ mprj.PS_Rx_inst3.LUT_inst1.i3 _0044_ _0092_ _0739_/VDD _0739_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1007_ _0269_ _0076_ _0138_ _0239_ _0349_ _0350_ _1007_/VDD _1007_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xuser_project_wrapper_127 io_out[20] user_project_wrapper_127/VDD user_project_wrapper_127/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_116 io_out[9] user_project_wrapper_116/VDD user_project_wrapper_116/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_138 io_out[31] user_project_wrapper_138/VDD user_project_wrapper_138/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_149 la_data_out[4] user_project_wrapper_149/VDD user_project_wrapper_149/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xoutput50 net50 wbs_dat_o[22] output50/VDD output50/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput61 net61 wbs_dat_o[3] output61/VDD output61/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xuser_project_wrapper_105 io_oeb[33] user_project_wrapper_105/VDD user_project_wrapper_105/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_0987_ mprj.PS_R1_inst1.LUT_inst14.I1 _0330_ _0987_/VDD _0987_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1272_ _0201_ _0586_ _0242_ _0602_ _1272_/VDD _1272_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1410_ _0025_ net68 mprj.PS_Rx_inst5.LUT_inst1.i4 _1410_/VDD _1410_/VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1341_ _0651_ _0012_ _1341_/VDD _1341_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0772_ _0111_ _0122_ _0123_ _0124_ _0772_/VDD _0772_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0841_ mprj.PS_R1_inst1.LUT_inst10.I0 _0189_ _0841_/VDD _0841_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0910_ mprj.PS_R1_inst1.LUT_inst7.I1 _0113_ _0129_ _0256_ _0910_/VDD _0910_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1186_ _0449_ _0157_ _0521_ _1186_/VDD _1186_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1324_ net24 _0094_ _0642_ _0643_ _1324_/VDD _1324_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1255_ _0449_ _0586_ _1255_/VDD _1255_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1040_ _0381_ _0382_ _1040_/VDD _1040_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1238_ _0154_ mprj.PS_Rx_inst5.LUT_inst1.i3 _0451_ _0570_ _1238_/VDD _1238_/VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1307_ _0586_ _0380_ _0632_ mprj.PS_Rx_inst8.LUT_inst1.i4 _0050_ _0633_ _1307_/VDD
+ _1307_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0755_ _0106_ _0107_ _0755_/VDD _0755_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_0824_ _0172_ _0173_ _0824_/VDD _0824_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_1169_ _0112_ _0449_ _0114_ _0505_ _1169_/VDD _1169_/VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_0686_ _0033_ _0038_ _0042_ _0043_ _0686_/VDD _0686_/VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_1023_ _0297_ _0076_ _0138_ mprj.PS_R1_inst1.LUT_inst12.I1 _0364_ _0365_ _1023_/VDD
+ _1023_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_0738_ _0069_ _0072_ _0091_ net61 _0738_/VDD _0738_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0807_ _0156_ _0157_ _0807_/VDD _0807_/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
Xuser_project_wrapper_90 io_oeb[18] user_project_wrapper_90/VDD user_project_wrapper_90/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1006_ mprj.PS_R1_inst1.LUT_inst12.I1 _0081_ _0099_ _0349_ _1006_/VDD _1006_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xuser_project_wrapper_128 io_out[21] user_project_wrapper_128/VDD user_project_wrapper_128/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_117 io_out[10] user_project_wrapper_117/VDD user_project_wrapper_117/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_139 io_out[32] user_project_wrapper_139/VDD user_project_wrapper_139/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xoutput51 net51 wbs_dat_o[23] output51/VDD output51/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput40 net40 wbs_dat_o[13] output40/VDD output40/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput62 net62 wbs_dat_o[4] output62/VDD output62/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xuser_project_wrapper_106 io_oeb[34] user_project_wrapper_106/VDD user_project_wrapper_106/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1340_ net17 _0270_ _0642_ _0651_ _1340_/VDD _1340_/VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1271_ _0187_ _0600_ _0331_ _0601_ _1271_/VDD _1271_/VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_0986_ mprj.PS_Rx_inst8.LUT_inst1.i3 _0044_ _0329_ _0986_/VDD _0986_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0840_ _0187_ _0068_ _0188_ _0840_/VDD _0840_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0771_ _0111_ _0122_ _0050_ _0123_ _0771_/VDD _0771_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1254_ _0451_ _0243_ _0585_ _1254_/VDD _1254_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1323_ _0636_ _0642_ _1323_/VDD _1323_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1185_ _0330_ _0149_ _0175_ _0520_ _1185_/VDD _1185_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0969_ _0280_ _0307_ _0312_ _0313_ _0969_/VDD _0969_/VSS gf180mcu_fd_sc_mcu7t5v0__xor3_4
X_1306_ _0322_ _0586_ _0631_ _0331_ _0632_ _1306_/VDD _1306_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_0823_ mprj.PS_Rx_inst4.LUT_inst1.i4 _0155_ _0172_ _0823_/VDD _0823_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_0685_ _0041_ _0032_ _0042_ _0685_/VDD _0685_/VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_0754_ mprj.PS_R1_inst1.LUT_inst5.I1 _0106_ _0754_/VDD _0754_/VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_1237_ _0270_ _0320_ _0337_ _0240_ _0568_ _0569_ _1237_/VDD _1237_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1168_ _0104_ _0450_ _0504_ _1168_/VDD _1168_/VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1099_ _0147_ _0248_ _0287_ _0127_ _0437_ _0438_ _1099_/VDD _1099_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1022_ mprj.PS_R1_inst1.LUT_inst13.I1 _0081_ _0099_ _0364_ _1022_/VDD _1022_/VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_0806_ _0154_ _0151_ _0155_ _0156_ _0806_/VDD _0806_/VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_0737_ _0067_ _0089_ _0090_ _0091_ _0737_/VDD _0737_/VSS gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xuser_project_wrapper_91 io_oeb[19] user_project_wrapper_91/VDD user_project_wrapper_91/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_80 io_oeb[8] user_project_wrapper_80/VDD user_project_wrapper_80/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
X_1005_ _0216_ _0115_ _0131_ _0189_ _0347_ _0348_ _1005_/VDD _1005_/VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xuser_project_wrapper_129 io_out[22] user_project_wrapper_129/VDD user_project_wrapper_129/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_project_wrapper_118 io_out[11] user_project_wrapper_118/VDD user_project_wrapper_118/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xoutput52 net52 wbs_dat_o[24] output52/VDD output52/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput41 net41 wbs_dat_o[14] output41/VDD output41/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xuser_project_wrapper_107 io_oeb[35] user_project_wrapper_107/VDD user_project_wrapper_107/VSS
+ gf180mcu_fd_sc_mcu7t5v0__tiel
Xoutput63 net63 wbs_dat_o[5] output63/VDD output63/VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
.ends

