VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_asic
  CLASS BLOCK ;
  FOREIGN user_proj_asic ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN A_PAD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 296.000 299.830 299.000 ;
    END
  END A_PAD
  PIN B_PAD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 1.000 145.270 4.000 ;
    END
  END B_PAD
  PIN OUT_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 146.240 299.000 146.840 ;
    END
  END OUT_1
  PIN OUT_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 153.040 4.000 153.640 ;
    END
  END OUT_2
  PIN sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END sel
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 296.000 6.810 299.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 294.640 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 294.640 181.510 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 288.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 294.640 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 294.640 184.810 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 296.000 154.930 299.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 1.000 293.390 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 0.070 6.500 299.850 288.560 ;
      LAYER met2 ;
        RECT 0.100 295.720 6.250 296.000 ;
        RECT 7.090 295.720 154.370 296.000 ;
        RECT 155.210 295.720 299.270 296.000 ;
        RECT 0.100 4.280 299.820 295.720 ;
        RECT 0.650 4.000 144.710 4.280 ;
        RECT 145.550 4.000 292.830 4.280 ;
        RECT 293.670 4.000 299.820 4.280 ;
      LAYER met3 ;
        RECT 4.000 154.040 296.000 288.485 ;
        RECT 4.400 152.640 296.000 154.040 ;
        RECT 4.000 147.240 296.000 152.640 ;
        RECT 4.000 145.840 295.600 147.240 ;
        RECT 4.000 10.715 296.000 145.840 ;
      LAYER met4 ;
        RECT 162.215 130.055 174.240 237.145 ;
        RECT 176.640 130.055 177.540 237.145 ;
        RECT 179.940 130.055 243.505 237.145 ;
  END
END user_proj_asic
END LIBRARY

