magic
tech sky130A
magscale 1 2
timestamp 1671619105
<< viali >>
rect 1593 57409 1627 57443
rect 2973 57409 3007 57443
rect 1777 57205 1811 57239
rect 2421 57205 2455 57239
rect 2145 56865 2179 56899
rect 2789 56865 2823 56899
rect 1961 56797 1995 56831
rect 58265 56797 58299 56831
rect 1593 56661 1627 56695
rect 2053 56661 2087 56695
rect 58173 56661 58207 56695
rect 58357 56457 58391 56491
rect 1685 56389 1719 56423
rect 1961 56117 1995 56151
rect 41797 48773 41831 48807
rect 36185 48705 36219 48739
rect 37657 48705 37691 48739
rect 38669 48705 38703 48739
rect 39681 48705 39715 48739
rect 40785 48705 40819 48739
rect 40969 48705 41003 48739
rect 42809 48705 42843 48739
rect 44005 48705 44039 48739
rect 36277 48637 36311 48671
rect 37565 48637 37599 48671
rect 38761 48637 38795 48671
rect 39589 48637 39623 48671
rect 42901 48637 42935 48671
rect 44097 48637 44131 48671
rect 35357 48569 35391 48603
rect 36553 48569 36587 48603
rect 39037 48569 39071 48603
rect 40049 48569 40083 48603
rect 33701 48501 33735 48535
rect 34253 48501 34287 48535
rect 34805 48501 34839 48535
rect 37933 48501 37967 48535
rect 43177 48501 43211 48535
rect 44373 48501 44407 48535
rect 35449 48229 35483 48263
rect 36461 48229 36495 48263
rect 40601 48229 40635 48263
rect 41613 48229 41647 48263
rect 33885 48161 33919 48195
rect 34161 48161 34195 48195
rect 34989 48161 35023 48195
rect 36001 48161 36035 48195
rect 40141 48161 40175 48195
rect 41153 48161 41187 48195
rect 33793 48093 33827 48127
rect 35081 48093 35115 48127
rect 36093 48093 36127 48127
rect 40233 48093 40267 48127
rect 41245 48093 41279 48127
rect 37013 48025 37047 48059
rect 37565 48025 37599 48059
rect 33149 47957 33183 47991
rect 38117 47957 38151 47991
rect 42073 47957 42107 47991
rect 39313 47753 39347 47787
rect 41337 47753 41371 47787
rect 34897 47685 34931 47719
rect 36645 47685 36679 47719
rect 32505 47617 32539 47651
rect 33517 47617 33551 47651
rect 35817 47617 35851 47651
rect 37657 47617 37691 47651
rect 38945 47617 38979 47651
rect 40969 47617 41003 47651
rect 42809 47617 42843 47651
rect 44281 47617 44315 47651
rect 44465 47617 44499 47651
rect 46489 47617 46523 47651
rect 32597 47549 32631 47583
rect 32873 47549 32907 47583
rect 33425 47549 33459 47583
rect 35725 47549 35759 47583
rect 37749 47549 37783 47583
rect 38853 47549 38887 47583
rect 40877 47549 40911 47583
rect 42901 47549 42935 47583
rect 45293 47549 45327 47583
rect 46397 47549 46431 47583
rect 33885 47481 33919 47515
rect 36185 47481 36219 47515
rect 38025 47481 38059 47515
rect 34621 47413 34655 47447
rect 39865 47413 39899 47447
rect 41889 47413 41923 47447
rect 43085 47413 43119 47447
rect 46857 47413 46891 47447
rect 36829 47209 36863 47243
rect 38025 47209 38059 47243
rect 34161 47141 34195 47175
rect 39313 47141 39347 47175
rect 42993 47141 43027 47175
rect 45753 47141 45787 47175
rect 46765 47141 46799 47175
rect 32045 47073 32079 47107
rect 34345 47073 34379 47107
rect 36645 47073 36679 47107
rect 37841 47073 37875 47107
rect 38853 47073 38887 47107
rect 40325 47073 40359 47107
rect 40785 47073 40819 47107
rect 42533 47073 42567 47107
rect 45293 47073 45327 47107
rect 46305 47073 46339 47107
rect 32229 47005 32263 47039
rect 32321 47005 32355 47039
rect 34069 47005 34103 47039
rect 34897 47005 34931 47039
rect 34990 47005 35024 47039
rect 35362 47005 35396 47039
rect 36093 47005 36127 47039
rect 36921 47005 36955 47039
rect 38117 47005 38151 47039
rect 38577 47005 38611 47039
rect 38669 47005 38703 47039
rect 40049 47005 40083 47039
rect 40141 47005 40175 47039
rect 40969 47005 41003 47039
rect 41061 47005 41095 47039
rect 42625 47005 42659 47039
rect 45385 47005 45419 47039
rect 46397 47005 46431 47039
rect 32873 46937 32907 46971
rect 33425 46937 33459 46971
rect 34345 46937 34379 46971
rect 35173 46937 35207 46971
rect 35265 46937 35299 46971
rect 36645 46937 36679 46971
rect 32045 46869 32079 46903
rect 35541 46869 35575 46903
rect 37841 46869 37875 46903
rect 38853 46869 38887 46903
rect 40325 46869 40359 46903
rect 40785 46869 40819 46903
rect 41613 46869 41647 46903
rect 43545 46869 43579 46903
rect 44005 46869 44039 46903
rect 44649 46869 44683 46903
rect 32597 46665 32631 46699
rect 34713 46665 34747 46699
rect 38117 46665 38151 46699
rect 39221 46665 39255 46699
rect 40325 46665 40359 46699
rect 41429 46665 41463 46699
rect 43269 46665 43303 46699
rect 44465 46665 44499 46699
rect 31217 46597 31251 46631
rect 40049 46597 40083 46631
rect 41061 46597 41095 46631
rect 42993 46597 43027 46631
rect 44097 46597 44131 46631
rect 46029 46597 46063 46631
rect 32321 46529 32355 46563
rect 33241 46529 33275 46563
rect 33609 46529 33643 46563
rect 34621 46529 34655 46563
rect 35541 46529 35575 46563
rect 36093 46529 36127 46563
rect 37473 46529 37507 46563
rect 37621 46529 37655 46563
rect 37749 46529 37783 46563
rect 37841 46529 37875 46563
rect 37979 46529 38013 46563
rect 38577 46529 38611 46563
rect 38670 46529 38704 46563
rect 38853 46529 38887 46563
rect 38945 46529 38979 46563
rect 39042 46529 39076 46563
rect 39681 46529 39715 46563
rect 39774 46529 39808 46563
rect 39957 46529 39991 46563
rect 40146 46529 40180 46563
rect 40785 46529 40819 46563
rect 40933 46529 40967 46563
rect 41153 46529 41187 46563
rect 41250 46529 41284 46563
rect 42625 46529 42659 46563
rect 42718 46529 42752 46563
rect 42901 46529 42935 46563
rect 43131 46529 43165 46563
rect 43821 46529 43855 46563
rect 43969 46529 44003 46563
rect 44189 46529 44223 46563
rect 44286 46529 44320 46563
rect 45017 46529 45051 46563
rect 45201 46529 45235 46563
rect 47869 46529 47903 46563
rect 48053 46529 48087 46563
rect 49341 46529 49375 46563
rect 33333 46461 33367 46495
rect 33517 46461 33551 46495
rect 35357 46461 35391 46495
rect 35909 46461 35943 46495
rect 48789 46461 48823 46495
rect 49525 46461 49559 46495
rect 31769 46325 31803 46359
rect 41889 46325 41923 46359
rect 31769 46121 31803 46155
rect 32965 46121 32999 46155
rect 33701 46121 33735 46155
rect 41061 46121 41095 46155
rect 41981 46121 42015 46155
rect 44281 46121 44315 46155
rect 47041 46053 47075 46087
rect 31033 45985 31067 46019
rect 36185 45985 36219 46019
rect 36461 45985 36495 46019
rect 37749 45985 37783 46019
rect 38577 45985 38611 46019
rect 42901 45985 42935 46019
rect 31493 45917 31527 45951
rect 31585 45917 31619 45951
rect 32321 45917 32355 45951
rect 32469 45917 32503 45951
rect 32786 45917 32820 45951
rect 33425 45917 33459 45951
rect 34161 45917 34195 45951
rect 35265 45917 35299 45951
rect 35817 45917 35851 45951
rect 36093 45917 36127 45951
rect 36737 45917 36771 45951
rect 37565 45917 37599 45951
rect 38393 45917 38427 45951
rect 38853 45917 38887 45951
rect 39221 45917 39255 45951
rect 40417 45917 40451 45951
rect 40510 45917 40544 45951
rect 40882 45917 40916 45951
rect 42625 45917 42659 45951
rect 43637 45917 43671 45951
rect 43785 45917 43819 45951
rect 44143 45917 44177 45951
rect 48513 45917 48547 45951
rect 48697 45917 48731 45951
rect 31769 45849 31803 45883
rect 32597 45849 32631 45883
rect 32689 45849 32723 45883
rect 33701 45849 33735 45883
rect 40693 45849 40727 45883
rect 40785 45849 40819 45883
rect 41705 45849 41739 45883
rect 43913 45849 43947 45883
rect 44005 45849 44039 45883
rect 46213 45849 46247 45883
rect 46857 45849 46891 45883
rect 33517 45781 33551 45815
rect 45293 45781 45327 45815
rect 49525 45781 49559 45815
rect 50445 45781 50479 45815
rect 51641 45781 51675 45815
rect 34253 45577 34287 45611
rect 41889 45577 41923 45611
rect 43453 45577 43487 45611
rect 44097 45577 44131 45611
rect 48329 45577 48363 45611
rect 36737 45509 36771 45543
rect 39865 45509 39899 45543
rect 40601 45509 40635 45543
rect 30573 45441 30607 45475
rect 31033 45441 31067 45475
rect 31217 45441 31251 45475
rect 31309 45441 31343 45475
rect 32413 45441 32447 45475
rect 32781 45441 32815 45475
rect 33333 45441 33367 45475
rect 34161 45441 34195 45475
rect 34437 45441 34471 45475
rect 35081 45441 35115 45475
rect 36645 45441 36679 45475
rect 36921 45441 36955 45475
rect 38209 45441 38243 45475
rect 39589 45441 39623 45475
rect 40325 45441 40359 45475
rect 40473 45441 40507 45475
rect 40693 45441 40727 45475
rect 40790 45441 40824 45475
rect 41797 45441 41831 45475
rect 42073 45441 42107 45475
rect 43177 45441 43211 45475
rect 43913 45441 43947 45475
rect 44189 45441 44223 45475
rect 45017 45441 45051 45475
rect 46305 45441 46339 45475
rect 47961 45441 47995 45475
rect 49341 45441 49375 45475
rect 50721 45441 50755 45475
rect 34989 45373 35023 45407
rect 38117 45373 38151 45407
rect 39865 45373 39899 45407
rect 43453 45373 43487 45407
rect 44925 45373 44959 45407
rect 46213 45373 46247 45407
rect 48053 45373 48087 45407
rect 49525 45373 49559 45407
rect 50905 45373 50939 45407
rect 51549 45373 51583 45407
rect 34437 45305 34471 45339
rect 36001 45305 36035 45339
rect 36921 45305 36955 45339
rect 39037 45305 39071 45339
rect 40969 45305 41003 45339
rect 42073 45305 42107 45339
rect 42717 45305 42751 45339
rect 43913 45305 43947 45339
rect 45385 45305 45419 45339
rect 52009 45305 52043 45339
rect 31033 45237 31067 45271
rect 35357 45237 35391 45271
rect 37473 45237 37507 45271
rect 38485 45237 38519 45271
rect 39681 45237 39715 45271
rect 43269 45237 43303 45271
rect 46581 45237 46615 45271
rect 34069 45033 34103 45067
rect 40049 45033 40083 45067
rect 40693 45033 40727 45067
rect 43821 45033 43855 45067
rect 47133 45033 47167 45067
rect 50905 45033 50939 45067
rect 42809 44965 42843 44999
rect 31861 44897 31895 44931
rect 35725 44897 35759 44931
rect 38025 44897 38059 44931
rect 38669 44897 38703 44931
rect 43361 44897 43395 44931
rect 46305 44897 46339 44931
rect 48513 44897 48547 44931
rect 50629 44897 50663 44931
rect 52009 44897 52043 44931
rect 52285 44897 52319 44931
rect 31125 44829 31159 44863
rect 31677 44829 31711 44863
rect 32045 44829 32079 44863
rect 32597 44829 32631 44863
rect 32781 44829 32815 44863
rect 33425 44829 33459 44863
rect 33518 44829 33552 44863
rect 33890 44829 33924 44863
rect 35909 44829 35943 44863
rect 37289 44829 37323 44863
rect 37841 44829 37875 44863
rect 38117 44829 38151 44863
rect 38761 44829 38795 44863
rect 41613 44829 41647 44863
rect 42165 44829 42199 44863
rect 42258 44829 42292 44863
rect 42441 44829 42475 44863
rect 42671 44829 42705 44863
rect 43453 44829 43487 44863
rect 45293 44829 45327 44863
rect 45477 44829 45511 44863
rect 48421 44829 48455 44863
rect 50537 44829 50571 44863
rect 51917 44829 51951 44863
rect 33701 44761 33735 44795
rect 33793 44761 33827 44795
rect 36645 44761 36679 44795
rect 42533 44761 42567 44795
rect 34897 44693 34931 44727
rect 41337 44693 41371 44727
rect 44373 44693 44407 44727
rect 47685 44693 47719 44727
rect 48789 44693 48823 44727
rect 49341 44693 49375 44727
rect 52929 44693 52963 44727
rect 32873 44489 32907 44523
rect 34437 44489 34471 44523
rect 36737 44489 36771 44523
rect 41429 44489 41463 44523
rect 42073 44489 42107 44523
rect 42809 44489 42843 44523
rect 47041 44489 47075 44523
rect 48421 44489 48455 44523
rect 36001 44421 36035 44455
rect 48145 44421 48179 44455
rect 49157 44421 49191 44455
rect 52101 44421 52135 44455
rect 31217 44353 31251 44387
rect 32597 44353 32631 44387
rect 33793 44353 33827 44387
rect 34989 44353 35023 44387
rect 35173 44353 35207 44387
rect 36645 44353 36679 44387
rect 36921 44353 36955 44387
rect 38209 44353 38243 44387
rect 38945 44353 38979 44387
rect 39129 44353 39163 44387
rect 40601 44353 40635 44387
rect 42625 44353 42659 44387
rect 42901 44353 42935 44387
rect 43637 44353 43671 44387
rect 46857 44353 46891 44387
rect 47133 44353 47167 44387
rect 47777 44353 47811 44387
rect 47870 44353 47904 44387
rect 48053 44353 48087 44387
rect 48283 44353 48317 44387
rect 48881 44353 48915 44387
rect 48974 44353 49008 44387
rect 49249 44353 49283 44387
rect 49346 44353 49380 44387
rect 50261 44353 50295 44387
rect 50445 44353 50479 44387
rect 50537 44353 50571 44387
rect 51733 44353 51767 44387
rect 51826 44353 51860 44387
rect 52009 44353 52043 44387
rect 52239 44353 52273 44387
rect 53021 44353 53055 44387
rect 53205 44353 53239 44387
rect 54585 44353 54619 44387
rect 54953 44353 54987 44387
rect 31125 44285 31159 44319
rect 32873 44285 32907 44319
rect 33517 44285 33551 44319
rect 37933 44285 37967 44319
rect 38117 44285 38151 44319
rect 39957 44285 39991 44319
rect 40693 44285 40727 44319
rect 43545 44285 43579 44319
rect 44005 44285 44039 44319
rect 54033 44285 54067 44319
rect 55597 44285 55631 44319
rect 31585 44217 31619 44251
rect 36921 44217 36955 44251
rect 42625 44217 42659 44251
rect 46857 44217 46891 44251
rect 52377 44217 52411 44251
rect 32689 44149 32723 44183
rect 38025 44149 38059 44183
rect 40969 44149 41003 44183
rect 49525 44149 49559 44183
rect 50261 44149 50295 44183
rect 51089 44149 51123 44183
rect 34161 43945 34195 43979
rect 41521 43945 41555 43979
rect 42809 43945 42843 43979
rect 46305 43945 46339 43979
rect 46857 43945 46891 43979
rect 50997 43945 51031 43979
rect 51641 43945 51675 43979
rect 54033 43945 54067 43979
rect 34897 43877 34931 43911
rect 35541 43877 35575 43911
rect 36461 43877 36495 43911
rect 45753 43877 45787 43911
rect 52469 43877 52503 43911
rect 32597 43809 32631 43843
rect 40693 43809 40727 43843
rect 41705 43809 41739 43843
rect 45293 43809 45327 43843
rect 49157 43809 49191 43843
rect 53573 43809 53607 43843
rect 56517 43809 56551 43843
rect 31677 43741 31711 43775
rect 32045 43741 32079 43775
rect 37105 43741 37139 43775
rect 38301 43741 38335 43775
rect 38394 43741 38428 43775
rect 38766 43741 38800 43775
rect 40601 43741 40635 43775
rect 41429 43741 41463 43775
rect 42165 43741 42199 43775
rect 42313 43741 42347 43775
rect 42441 43741 42475 43775
rect 42671 43741 42705 43775
rect 43269 43741 43303 43775
rect 45385 43741 45419 43775
rect 47036 43741 47070 43775
rect 47408 43741 47442 43775
rect 47501 43741 47535 43775
rect 49249 43741 49283 43775
rect 50353 43741 50387 43775
rect 50501 43741 50535 43775
rect 50818 43741 50852 43775
rect 51641 43741 51675 43775
rect 51917 43741 51951 43775
rect 53665 43741 53699 43775
rect 55597 43741 55631 43775
rect 55781 43741 55815 43775
rect 33241 43673 33275 43707
rect 36185 43673 36219 43707
rect 37473 43673 37507 43707
rect 38577 43673 38611 43707
rect 38669 43673 38703 43707
rect 42533 43673 42567 43707
rect 44097 43673 44131 43707
rect 47133 43673 47167 43707
rect 47225 43673 47259 43707
rect 48237 43673 48271 43707
rect 50629 43673 50663 43707
rect 50721 43673 50755 43707
rect 33517 43605 33551 43639
rect 38945 43605 38979 43639
rect 39405 43605 39439 43639
rect 40969 43605 41003 43639
rect 41705 43605 41739 43639
rect 43453 43605 43487 43639
rect 44557 43605 44591 43639
rect 48329 43605 48363 43639
rect 49617 43605 49651 43639
rect 51825 43605 51859 43639
rect 52929 43605 52963 43639
rect 54493 43605 54527 43639
rect 34345 43401 34379 43435
rect 36277 43401 36311 43435
rect 38577 43401 38611 43435
rect 40601 43401 40635 43435
rect 41797 43401 41831 43435
rect 43269 43401 43303 43435
rect 44373 43401 44407 43435
rect 46305 43401 46339 43435
rect 47133 43401 47167 43435
rect 48145 43401 48179 43435
rect 54033 43401 54067 43435
rect 36553 43333 36587 43367
rect 39497 43333 39531 43367
rect 41984 43333 42018 43367
rect 42901 43333 42935 43367
rect 44005 43333 44039 43367
rect 44097 43333 44131 43367
rect 30757 43265 30791 43299
rect 32965 43265 32999 43299
rect 33977 43265 34011 43299
rect 34989 43265 35023 43299
rect 35082 43265 35116 43299
rect 35265 43265 35299 43299
rect 35357 43265 35391 43299
rect 35493 43265 35527 43299
rect 36415 43265 36449 43299
rect 36645 43265 36679 43299
rect 36773 43265 36807 43299
rect 36921 43265 36955 43299
rect 37749 43265 37783 43299
rect 39222 43265 39256 43299
rect 39957 43265 39991 43299
rect 40050 43265 40084 43299
rect 40233 43265 40267 43299
rect 40325 43265 40359 43299
rect 40463 43265 40497 43299
rect 41705 43265 41739 43299
rect 42625 43265 42659 43299
rect 42718 43265 42752 43299
rect 42993 43265 43027 43299
rect 43090 43265 43124 43299
rect 43729 43265 43763 43299
rect 43877 43265 43911 43299
rect 44194 43265 44228 43299
rect 45017 43265 45051 43299
rect 46857 43265 46891 43299
rect 48053 43265 48087 43299
rect 48329 43265 48363 43299
rect 48789 43265 48823 43299
rect 50077 43265 50111 43299
rect 51549 43265 51583 43299
rect 54953 43265 54987 43299
rect 30665 43197 30699 43231
rect 31125 43197 31159 43231
rect 32873 43197 32907 43231
rect 33885 43197 33919 43231
rect 37657 43197 37691 43231
rect 39497 43197 39531 43231
rect 44925 43197 44959 43231
rect 47133 43197 47167 43231
rect 49985 43197 50019 43231
rect 51273 43197 51307 43231
rect 52101 43197 52135 43231
rect 55045 43197 55079 43231
rect 55321 43197 55355 43231
rect 33333 43129 33367 43163
rect 41981 43129 42015 43163
rect 45385 43129 45419 43163
rect 48329 43129 48363 43163
rect 50445 43129 50479 43163
rect 35633 43061 35667 43095
rect 39313 43061 39347 43095
rect 41153 43061 41187 43095
rect 46949 43061 46983 43095
rect 48973 43061 49007 43095
rect 52929 43061 52963 43095
rect 53481 43061 53515 43095
rect 55781 43061 55815 43095
rect 31125 42857 31159 42891
rect 33241 42857 33275 42891
rect 37013 42857 37047 42891
rect 37105 42857 37139 42891
rect 42901 42857 42935 42891
rect 44373 42857 44407 42891
rect 48513 42857 48547 42891
rect 48605 42857 48639 42891
rect 49801 42857 49835 42891
rect 53757 42857 53791 42891
rect 54861 42857 54895 42891
rect 32689 42789 32723 42823
rect 34161 42789 34195 42823
rect 36369 42789 36403 42823
rect 38577 42789 38611 42823
rect 52377 42789 52411 42823
rect 56425 42789 56459 42823
rect 30757 42721 30791 42755
rect 34345 42721 34379 42755
rect 36921 42721 36955 42755
rect 38117 42721 38151 42755
rect 44189 42721 44223 42755
rect 48697 42721 48731 42755
rect 51917 42721 51951 42755
rect 55965 42721 55999 42755
rect 57161 42721 57195 42755
rect 30849 42653 30883 42687
rect 32045 42653 32079 42687
rect 32138 42653 32172 42687
rect 32413 42653 32447 42687
rect 32510 42653 32544 42687
rect 34069 42653 34103 42687
rect 35081 42653 35115 42687
rect 35174 42653 35208 42687
rect 35546 42653 35580 42687
rect 36185 42653 36219 42687
rect 37197 42653 37231 42687
rect 38209 42653 38243 42687
rect 41981 42653 42015 42687
rect 42717 42653 42751 42687
rect 43453 42653 43487 42687
rect 43729 42653 43763 42687
rect 44465 42653 44499 42687
rect 45753 42653 45787 42687
rect 45937 42653 45971 42687
rect 48421 42653 48455 42687
rect 49157 42653 49191 42687
rect 49250 42653 49284 42687
rect 49433 42653 49467 42687
rect 49663 42653 49697 42687
rect 52009 42653 52043 42687
rect 53113 42653 53147 42687
rect 53206 42653 53240 42687
rect 53481 42653 53515 42687
rect 53619 42653 53653 42687
rect 54217 42653 54251 42687
rect 54401 42653 54435 42687
rect 54493 42653 54527 42687
rect 54585 42653 54619 42687
rect 56057 42653 56091 42687
rect 57253 42653 57287 42687
rect 32321 42585 32355 42619
rect 34345 42585 34379 42619
rect 35357 42585 35391 42619
rect 35449 42585 35483 42619
rect 44189 42585 44223 42619
rect 46765 42585 46799 42619
rect 47685 42585 47719 42619
rect 49525 42585 49559 42619
rect 50353 42585 50387 42619
rect 50905 42585 50939 42619
rect 53389 42585 53423 42619
rect 35725 42517 35759 42551
rect 39037 42517 39071 42551
rect 40049 42517 40083 42551
rect 42165 42517 42199 42551
rect 43551 42517 43585 42551
rect 43637 42517 43671 42551
rect 58081 42517 58115 42551
rect 31769 42313 31803 42347
rect 32505 42313 32539 42347
rect 34897 42313 34931 42347
rect 36553 42313 36587 42347
rect 39773 42313 39807 42347
rect 44005 42313 44039 42347
rect 45569 42313 45603 42347
rect 47133 42313 47167 42347
rect 50261 42313 50295 42347
rect 53205 42313 53239 42347
rect 54769 42313 54803 42347
rect 55781 42313 55815 42347
rect 42073 42245 42107 42279
rect 43729 42245 43763 42279
rect 48145 42245 48179 42279
rect 55229 42245 55263 42279
rect 56333 42245 56367 42279
rect 29837 42177 29871 42211
rect 31493 42177 31527 42211
rect 32413 42177 32447 42211
rect 34621 42177 34655 42211
rect 34713 42177 34747 42211
rect 35725 42177 35759 42211
rect 36277 42177 36311 42211
rect 37473 42177 37507 42211
rect 38945 42177 38979 42211
rect 40601 42177 40635 42211
rect 41797 42177 41831 42211
rect 41889 42177 41923 42211
rect 43361 42177 43395 42211
rect 43454 42177 43488 42211
rect 43637 42177 43671 42211
rect 43867 42177 43901 42211
rect 45201 42177 45235 42211
rect 46949 42177 46983 42211
rect 47225 42177 47259 42211
rect 47956 42177 47990 42211
rect 48053 42177 48087 42211
rect 48273 42177 48307 42211
rect 48421 42177 48455 42211
rect 49065 42177 49099 42211
rect 49249 42177 49283 42211
rect 49341 42177 49375 42211
rect 49433 42177 49467 42211
rect 50905 42177 50939 42211
rect 52929 42177 52963 42211
rect 53021 42177 53055 42211
rect 54125 42177 54159 42211
rect 54273 42177 54307 42211
rect 54401 42177 54435 42211
rect 54493 42177 54527 42211
rect 54590 42177 54624 42211
rect 29745 42109 29779 42143
rect 30205 42109 30239 42143
rect 31769 42109 31803 42143
rect 34897 42109 34931 42143
rect 38853 42109 38887 42143
rect 40509 42109 40543 42143
rect 42809 42109 42843 42143
rect 45109 42109 45143 42143
rect 50997 42109 51031 42143
rect 51273 42109 51307 42143
rect 52285 42109 52319 42143
rect 53205 42109 53239 42143
rect 39313 42041 39347 42075
rect 40969 42041 41003 42075
rect 46949 42041 46983 42075
rect 31585 41973 31619 42007
rect 34161 41973 34195 42007
rect 37657 41973 37691 42007
rect 38209 41973 38243 42007
rect 42073 41973 42107 42007
rect 44465 41973 44499 42007
rect 47777 41973 47811 42007
rect 49709 41973 49743 42007
rect 51825 41973 51859 42007
rect 33701 41769 33735 41803
rect 36645 41769 36679 41803
rect 40785 41769 40819 41803
rect 48605 41769 48639 41803
rect 49157 41769 49191 41803
rect 54677 41769 54711 41803
rect 31033 41701 31067 41735
rect 42993 41701 43027 41735
rect 52745 41701 52779 41735
rect 28917 41633 28951 41667
rect 29193 41633 29227 41667
rect 30021 41633 30055 41667
rect 31861 41633 31895 41667
rect 33333 41633 33367 41667
rect 36001 41633 36035 41667
rect 38025 41633 38059 41667
rect 38669 41633 38703 41667
rect 43913 41633 43947 41667
rect 44189 41633 44223 41667
rect 45385 41633 45419 41667
rect 46305 41633 46339 41667
rect 47501 41633 47535 41667
rect 50445 41633 50479 41667
rect 53205 41633 53239 41667
rect 54033 41633 54067 41667
rect 56149 41633 56183 41667
rect 57069 41633 57103 41667
rect 28825 41565 28859 41599
rect 30113 41565 30147 41599
rect 30941 41565 30975 41599
rect 31769 41565 31803 41599
rect 32229 41565 32263 41599
rect 32781 41565 32815 41599
rect 33425 41565 33459 41599
rect 34989 41565 35023 41599
rect 35173 41565 35207 41599
rect 36461 41565 36495 41599
rect 37473 41565 37507 41599
rect 37841 41565 37875 41599
rect 38117 41565 38151 41599
rect 38761 41565 38795 41599
rect 40141 41565 40175 41599
rect 40261 41565 40295 41599
rect 40506 41565 40540 41599
rect 40645 41565 40679 41599
rect 41337 41565 41371 41599
rect 42349 41565 42383 41599
rect 42442 41565 42476 41599
rect 42625 41565 42659 41599
rect 42814 41565 42848 41599
rect 43821 41565 43855 41599
rect 45477 41565 45511 41599
rect 47409 41565 47443 41599
rect 48329 41565 48363 41599
rect 49530 41565 49564 41599
rect 50537 41565 50571 41599
rect 52101 41565 52135 41599
rect 52194 41565 52228 41599
rect 52469 41565 52503 41599
rect 52566 41565 52600 41599
rect 53757 41565 53791 41599
rect 53941 41565 53975 41599
rect 54130 41565 54164 41599
rect 56241 41565 56275 41599
rect 40417 41497 40451 41531
rect 41705 41497 41739 41531
rect 42717 41497 42751 41531
rect 49157 41497 49191 41531
rect 49341 41497 49375 41531
rect 49433 41497 49467 41531
rect 52377 41497 52411 41531
rect 54033 41497 54067 41531
rect 30481 41429 30515 41463
rect 47777 41429 47811 41463
rect 50905 41429 50939 41463
rect 51365 41429 51399 41463
rect 32873 41225 32907 41259
rect 33885 41225 33919 41259
rect 36553 41225 36587 41259
rect 38853 41225 38887 41259
rect 40693 41225 40727 41259
rect 47869 41225 47903 41259
rect 49249 41225 49283 41259
rect 50905 41225 50939 41259
rect 55597 41225 55631 41259
rect 35633 41157 35667 41191
rect 38485 41157 38519 41191
rect 41889 41157 41923 41191
rect 42993 41157 43027 41191
rect 47225 41157 47259 41191
rect 51733 41157 51767 41191
rect 53021 41157 53055 41191
rect 32505 41089 32539 41123
rect 33517 41089 33551 41123
rect 35444 41089 35478 41123
rect 35541 41089 35575 41123
rect 35816 41089 35850 41123
rect 35909 41089 35943 41123
rect 36369 41089 36403 41123
rect 37473 41089 37507 41123
rect 37565 41089 37599 41123
rect 37749 41089 37783 41123
rect 38209 41089 38243 41123
rect 38347 41089 38381 41123
rect 38606 41089 38640 41123
rect 38715 41089 38749 41123
rect 39865 41089 39899 41123
rect 41797 41089 41831 41123
rect 42073 41089 42107 41123
rect 42625 41089 42659 41123
rect 42718 41089 42752 41123
rect 42901 41089 42935 41123
rect 43131 41089 43165 41123
rect 43913 41089 43947 41123
rect 46581 41089 46615 41123
rect 48513 41089 48547 41123
rect 50813 41089 50847 41123
rect 51089 41089 51123 41123
rect 51549 41089 51583 41123
rect 51821 41089 51855 41123
rect 52285 41089 52319 41123
rect 53849 41089 53883 41123
rect 55229 41089 55263 41123
rect 32413 41021 32447 41055
rect 33609 41021 33643 41055
rect 40141 41021 40175 41055
rect 43821 41021 43855 41055
rect 44281 41021 44315 41055
rect 46305 41021 46339 41055
rect 48789 41021 48823 41055
rect 50261 41021 50295 41055
rect 55137 41021 55171 41055
rect 35265 40953 35299 40987
rect 37749 40953 37783 40987
rect 42073 40953 42107 40987
rect 43269 40953 43303 40987
rect 48605 40953 48639 40987
rect 39313 40885 39347 40919
rect 39957 40885 39991 40919
rect 40049 40885 40083 40919
rect 48697 40885 48731 40919
rect 51089 40885 51123 40919
rect 51549 40885 51583 40919
rect 53113 40885 53147 40919
rect 54033 40885 54067 40919
rect 56057 40885 56091 40919
rect 56609 40885 56643 40919
rect 29101 40681 29135 40715
rect 31217 40681 31251 40715
rect 32321 40681 32355 40715
rect 35173 40681 35207 40715
rect 35265 40681 35299 40715
rect 36277 40681 36311 40715
rect 36921 40681 36955 40715
rect 37933 40681 37967 40715
rect 38669 40681 38703 40715
rect 40141 40681 40175 40715
rect 53389 40681 53423 40715
rect 42625 40613 42659 40647
rect 45753 40613 45787 40647
rect 52653 40613 52687 40647
rect 28733 40545 28767 40579
rect 32965 40545 32999 40579
rect 35357 40545 35391 40579
rect 37105 40545 37139 40579
rect 37841 40545 37875 40579
rect 45293 40545 45327 40579
rect 46581 40545 46615 40579
rect 50905 40545 50939 40579
rect 53481 40545 53515 40579
rect 28825 40477 28859 40511
rect 30573 40477 30607 40511
rect 30666 40477 30700 40511
rect 31079 40477 31113 40511
rect 32505 40477 32539 40511
rect 33149 40477 33183 40511
rect 33241 40477 33275 40511
rect 35081 40477 35115 40511
rect 36829 40477 36863 40511
rect 38025 40477 38059 40511
rect 38117 40477 38151 40511
rect 40693 40477 40727 40511
rect 42349 40477 42383 40511
rect 45385 40477 45419 40511
rect 46673 40477 46707 40511
rect 48508 40477 48542 40511
rect 48605 40477 48639 40511
rect 48825 40477 48859 40511
rect 48973 40477 49007 40511
rect 50629 40477 50663 40511
rect 52009 40477 52043 40511
rect 52102 40477 52136 40511
rect 52377 40477 52411 40511
rect 52474 40477 52508 40511
rect 53205 40477 53239 40511
rect 53297 40477 53331 40511
rect 53941 40477 53975 40511
rect 54034 40477 54068 40511
rect 54217 40477 54251 40511
rect 54406 40477 54440 40511
rect 55597 40477 55631 40511
rect 57253 40477 57287 40511
rect 57437 40477 57471 40511
rect 30849 40409 30883 40443
rect 30941 40409 30975 40443
rect 42625 40409 42659 40443
rect 48697 40409 48731 40443
rect 52285 40409 52319 40443
rect 54309 40409 54343 40443
rect 56609 40409 56643 40443
rect 32965 40341 32999 40375
rect 37105 40341 37139 40375
rect 39221 40341 39255 40375
rect 40785 40341 40819 40375
rect 42441 40341 42475 40375
rect 47501 40341 47535 40375
rect 48329 40341 48363 40375
rect 49709 40341 49743 40375
rect 51457 40341 51491 40375
rect 54585 40341 54619 40375
rect 58265 40341 58299 40375
rect 41882 40137 41916 40171
rect 43269 40137 43303 40171
rect 44281 40137 44315 40171
rect 54033 40137 54067 40171
rect 57161 40137 57195 40171
rect 30297 40069 30331 40103
rect 31033 40069 31067 40103
rect 32597 40069 32631 40103
rect 32689 40069 32723 40103
rect 37749 40069 37783 40103
rect 41797 40069 41831 40103
rect 41981 40069 42015 40103
rect 42901 40069 42935 40103
rect 50997 40069 51031 40103
rect 30021 40001 30055 40035
rect 30757 40001 30791 40035
rect 30905 40001 30939 40035
rect 31125 40001 31159 40035
rect 31263 40001 31297 40035
rect 32500 40001 32534 40035
rect 32872 40001 32906 40035
rect 32965 40001 32999 40035
rect 33609 40001 33643 40035
rect 36093 40001 36127 40035
rect 37462 40001 37496 40035
rect 37621 40001 37655 40035
rect 37841 40001 37875 40035
rect 37979 40001 38013 40035
rect 38945 40001 38979 40035
rect 39865 40001 39899 40035
rect 41705 40001 41739 40035
rect 42625 40001 42659 40035
rect 42718 40001 42752 40035
rect 42993 40001 43027 40035
rect 43131 40001 43165 40035
rect 43913 40001 43947 40035
rect 46765 40001 46799 40035
rect 48605 40001 48639 40035
rect 49617 40001 49651 40035
rect 51917 40001 51951 40035
rect 53021 40001 53055 40035
rect 53757 40001 53791 40035
rect 54953 40001 54987 40035
rect 56793 40001 56827 40035
rect 30297 39933 30331 39967
rect 33517 39933 33551 39967
rect 35909 39933 35943 39967
rect 36829 39933 36863 39967
rect 43821 39933 43855 39967
rect 48513 39933 48547 39967
rect 49525 39933 49559 39967
rect 51273 39933 51307 39967
rect 54033 39933 54067 39967
rect 54861 39933 54895 39967
rect 56701 39933 56735 39967
rect 31401 39865 31435 39899
rect 32321 39865 32355 39899
rect 33977 39865 34011 39899
rect 40785 39865 40819 39899
rect 48973 39865 49007 39899
rect 49985 39865 50019 39899
rect 53205 39865 53239 39899
rect 55321 39865 55355 39899
rect 30113 39797 30147 39831
rect 38117 39797 38151 39831
rect 47777 39797 47811 39831
rect 53849 39797 53883 39831
rect 55781 39797 55815 39831
rect 29009 39593 29043 39627
rect 31677 39593 31711 39627
rect 32597 39593 32631 39627
rect 34069 39593 34103 39627
rect 36093 39593 36127 39627
rect 37013 39593 37047 39627
rect 29101 39525 29135 39559
rect 39497 39525 39531 39559
rect 43361 39525 43395 39559
rect 44649 39525 44683 39559
rect 47225 39525 47259 39559
rect 48697 39525 48731 39559
rect 53481 39525 53515 39559
rect 29193 39457 29227 39491
rect 33885 39457 33919 39491
rect 36829 39457 36863 39491
rect 38117 39457 38151 39491
rect 38853 39457 38887 39491
rect 44189 39457 44223 39491
rect 45569 39457 45603 39491
rect 46489 39457 46523 39491
rect 50353 39457 50387 39491
rect 52561 39457 52595 39491
rect 53389 39457 53423 39491
rect 53573 39457 53607 39491
rect 55689 39457 55723 39491
rect 28917 39389 28951 39423
rect 29837 39389 29871 39423
rect 30849 39389 30883 39423
rect 33793 39389 33827 39423
rect 35449 39389 35483 39423
rect 35542 39389 35576 39423
rect 35817 39389 35851 39423
rect 35955 39389 35989 39423
rect 37105 39389 37139 39423
rect 38025 39389 38059 39423
rect 39313 39389 39347 39423
rect 39497 39389 39531 39423
rect 40141 39389 40175 39423
rect 41792 39389 41826 39423
rect 41981 39389 42015 39423
rect 42109 39389 42143 39423
rect 42268 39389 42302 39423
rect 42717 39389 42751 39423
rect 42837 39389 42871 39423
rect 43085 39389 43119 39423
rect 43182 39389 43216 39423
rect 44281 39389 44315 39423
rect 45661 39389 45695 39423
rect 46949 39389 46983 39423
rect 47041 39389 47075 39423
rect 48053 39389 48087 39423
rect 48201 39389 48235 39423
rect 48518 39389 48552 39423
rect 51917 39389 51951 39423
rect 53297 39389 53331 39423
rect 54033 39389 54067 39423
rect 54126 39389 54160 39423
rect 54309 39389 54343 39423
rect 54539 39389 54573 39423
rect 55781 39389 55815 39423
rect 57069 39389 57103 39423
rect 57253 39389 57287 39423
rect 31401 39321 31435 39355
rect 32321 39321 32355 39355
rect 35725 39321 35759 39355
rect 41153 39321 41187 39355
rect 41889 39321 41923 39355
rect 42993 39321 43027 39355
rect 47225 39321 47259 39355
rect 48329 39321 48363 39355
rect 48421 39321 48455 39355
rect 49709 39321 49743 39355
rect 51641 39321 51675 39355
rect 54401 39321 54435 39355
rect 36829 39253 36863 39287
rect 41613 39253 41647 39287
rect 49157 39253 49191 39287
rect 51089 39253 51123 39287
rect 51739 39253 51773 39287
rect 51825 39253 51859 39287
rect 54677 39253 54711 39287
rect 56149 39253 56183 39287
rect 58081 39253 58115 39287
rect 30573 39049 30607 39083
rect 31585 39049 31619 39083
rect 32873 39049 32907 39083
rect 34437 39049 34471 39083
rect 35541 39049 35575 39083
rect 41981 39049 42015 39083
rect 46305 39049 46339 39083
rect 47133 39049 47167 39083
rect 48973 39049 49007 39083
rect 56885 39049 56919 39083
rect 36553 38981 36587 39015
rect 45109 38981 45143 39015
rect 48605 38981 48639 39015
rect 50261 38981 50295 39015
rect 54493 38981 54527 39015
rect 29745 38913 29779 38947
rect 30757 38913 30791 38947
rect 31493 38913 31527 38947
rect 31769 38913 31803 38947
rect 32965 38913 32999 38947
rect 34069 38913 34103 38947
rect 35265 38913 35299 38947
rect 36415 38913 36449 38947
rect 36645 38913 36679 38947
rect 36828 38913 36862 38947
rect 36921 38913 36955 38947
rect 38577 38913 38611 38947
rect 39221 38913 39255 38947
rect 41153 38913 41187 38947
rect 42625 38913 42659 38947
rect 42718 38913 42752 38947
rect 42901 38913 42935 38947
rect 42993 38913 43027 38947
rect 43131 38913 43165 38947
rect 44189 38913 44223 38947
rect 45017 38913 45051 38947
rect 45201 38913 45235 38947
rect 46489 38913 46523 38947
rect 46949 38913 46983 38947
rect 48329 38913 48363 38947
rect 48422 38913 48456 38947
rect 48697 38913 48731 38947
rect 48794 38913 48828 38947
rect 49985 38913 50019 38947
rect 50077 38913 50111 38947
rect 51089 38913 51123 38947
rect 53067 38913 53101 38947
rect 53205 38913 53239 38947
rect 53297 38913 53331 38947
rect 53480 38913 53514 38947
rect 53573 38913 53607 38947
rect 54217 38913 54251 38947
rect 54310 38913 54344 38947
rect 54585 38913 54619 38947
rect 54682 38913 54716 38947
rect 56517 38913 56551 38947
rect 30021 38845 30055 38879
rect 33977 38845 34011 38879
rect 35357 38845 35391 38879
rect 35541 38845 35575 38879
rect 39865 38845 39899 38879
rect 41061 38845 41095 38879
rect 44097 38845 44131 38879
rect 51181 38845 51215 38879
rect 51917 38845 51951 38879
rect 55321 38845 55355 38879
rect 56425 38845 56459 38879
rect 29837 38777 29871 38811
rect 43269 38777 43303 38811
rect 44557 38777 44591 38811
rect 57345 38777 57379 38811
rect 29929 38709 29963 38743
rect 31769 38709 31803 38743
rect 36277 38709 36311 38743
rect 37565 38709 37599 38743
rect 45661 38709 45695 38743
rect 47869 38709 47903 38743
rect 49433 38709 49467 38743
rect 50261 38709 50295 38743
rect 52929 38709 52963 38743
rect 54861 38709 54895 38743
rect 31309 38505 31343 38539
rect 33885 38505 33919 38539
rect 35357 38505 35391 38539
rect 35909 38505 35943 38539
rect 41061 38505 41095 38539
rect 47225 38505 47259 38539
rect 48145 38505 48179 38539
rect 50997 38505 51031 38539
rect 52009 38505 52043 38539
rect 53941 38505 53975 38539
rect 54033 38505 54067 38539
rect 56517 38505 56551 38539
rect 29009 38437 29043 38471
rect 32873 38437 32907 38471
rect 43913 38437 43947 38471
rect 49709 38437 49743 38471
rect 54585 38437 54619 38471
rect 33425 38369 33459 38403
rect 38577 38369 38611 38403
rect 43453 38369 43487 38403
rect 45753 38369 45787 38403
rect 46397 38369 46431 38403
rect 49249 38369 49283 38403
rect 52837 38369 52871 38403
rect 54125 38369 54159 38403
rect 55597 38369 55631 38403
rect 29193 38301 29227 38335
rect 30665 38301 30699 38335
rect 30813 38301 30847 38335
rect 31033 38301 31067 38335
rect 31171 38301 31205 38335
rect 32229 38301 32263 38335
rect 32322 38301 32356 38335
rect 32505 38301 32539 38335
rect 32694 38301 32728 38335
rect 33517 38301 33551 38335
rect 34897 38301 34931 38335
rect 35081 38301 35115 38335
rect 35909 38301 35943 38335
rect 36001 38301 36035 38335
rect 36645 38301 36679 38335
rect 36829 38301 36863 38335
rect 37565 38301 37599 38335
rect 37933 38301 37967 38335
rect 39129 38301 39163 38335
rect 39313 38301 39347 38335
rect 40417 38301 40451 38335
rect 40510 38301 40544 38335
rect 40693 38301 40727 38335
rect 40923 38301 40957 38335
rect 43545 38301 43579 38335
rect 45569 38301 45603 38335
rect 47409 38301 47443 38335
rect 47869 38301 47903 38335
rect 49341 38301 49375 38335
rect 50353 38301 50387 38335
rect 50446 38301 50480 38335
rect 50818 38301 50852 38335
rect 52745 38301 52779 38335
rect 53849 38301 53883 38335
rect 55689 38301 55723 38335
rect 29837 38233 29871 38267
rect 30941 38233 30975 38267
rect 32597 38233 32631 38267
rect 35449 38233 35483 38267
rect 36185 38233 36219 38267
rect 40785 38233 40819 38267
rect 41889 38233 41923 38267
rect 42533 38233 42567 38267
rect 42901 38233 42935 38267
rect 48145 38233 48179 38267
rect 50629 38233 50663 38267
rect 50721 38233 50755 38267
rect 51457 38233 51491 38267
rect 30113 38165 30147 38199
rect 36737 38165 36771 38199
rect 39497 38165 39531 38199
rect 41797 38165 41831 38199
rect 47961 38165 47995 38199
rect 48697 38165 48731 38199
rect 53113 38165 53147 38199
rect 56057 38165 56091 38199
rect 29285 37961 29319 37995
rect 31677 37961 31711 37995
rect 32781 37961 32815 37995
rect 33425 37961 33459 37995
rect 34437 37961 34471 37995
rect 39773 37961 39807 37995
rect 52285 37961 52319 37995
rect 54493 37961 54527 37995
rect 55045 37961 55079 37995
rect 32505 37893 32539 37927
rect 33577 37893 33611 37927
rect 33793 37893 33827 37927
rect 36001 37893 36035 37927
rect 40325 37893 40359 37927
rect 42901 37893 42935 37927
rect 42993 37893 43027 37927
rect 43821 37893 43855 37927
rect 47041 37893 47075 37927
rect 48513 37893 48547 37927
rect 49249 37893 49283 37927
rect 54033 37893 54067 37927
rect 29193 37825 29227 37859
rect 30113 37825 30147 37859
rect 30481 37825 30515 37859
rect 30941 37825 30975 37859
rect 31493 37825 31527 37859
rect 34621 37825 34655 37859
rect 34805 37825 34839 37859
rect 34897 37825 34931 37859
rect 35357 37825 35391 37859
rect 35633 37825 35667 37859
rect 36461 37825 36495 37859
rect 36645 37825 36679 37859
rect 37473 37825 37507 37859
rect 37657 37825 37691 37859
rect 37933 37825 37967 37859
rect 39497 37825 39531 37859
rect 39589 37825 39623 37859
rect 41245 37825 41279 37859
rect 42625 37825 42659 37859
rect 42718 37825 42752 37859
rect 43090 37825 43124 37859
rect 44833 37825 44867 37859
rect 46305 37825 46339 37859
rect 46489 37825 46523 37859
rect 46949 37825 46983 37859
rect 47225 37825 47259 37859
rect 48145 37825 48179 37859
rect 48238 37825 48272 37859
rect 48421 37825 48455 37859
rect 48610 37825 48644 37859
rect 50905 37825 50939 37859
rect 53205 37825 53239 37859
rect 55965 37825 55999 37859
rect 56977 37825 57011 37859
rect 30205 37757 30239 37791
rect 35817 37757 35851 37791
rect 36553 37757 36587 37791
rect 39773 37757 39807 37791
rect 44741 37757 44775 37791
rect 45661 37757 45695 37791
rect 50813 37757 50847 37791
rect 51273 37757 51307 37791
rect 53113 37757 53147 37791
rect 55873 37757 55907 37791
rect 56885 37757 56919 37791
rect 38117 37689 38151 37723
rect 47225 37689 47259 37723
rect 48789 37689 48823 37723
rect 56333 37689 56367 37723
rect 28733 37621 28767 37655
rect 33609 37621 33643 37655
rect 38669 37621 38703 37655
rect 40601 37621 40635 37655
rect 41521 37621 41555 37655
rect 43269 37621 43303 37655
rect 46489 37621 46523 37655
rect 49801 37621 49835 37655
rect 57253 37621 57287 37655
rect 29193 37417 29227 37451
rect 32321 37417 32355 37451
rect 34897 37417 34931 37451
rect 37381 37417 37415 37451
rect 41521 37417 41555 37451
rect 43729 37417 43763 37451
rect 46581 37417 46615 37451
rect 53481 37417 53515 37451
rect 56333 37417 56367 37451
rect 28457 37349 28491 37383
rect 33425 37349 33459 37383
rect 34253 37349 34287 37383
rect 35633 37349 35667 37383
rect 39497 37349 39531 37383
rect 40417 37349 40451 37383
rect 47777 37349 47811 37383
rect 30757 37281 30791 37315
rect 30941 37281 30975 37315
rect 32781 37281 32815 37315
rect 38209 37281 38243 37315
rect 38485 37281 38519 37315
rect 39037 37281 39071 37315
rect 43361 37281 43395 37315
rect 49433 37281 49467 37315
rect 51733 37281 51767 37315
rect 53665 37281 53699 37315
rect 55965 37281 55999 37315
rect 28181 37213 28215 37247
rect 28917 37213 28951 37247
rect 29009 37213 29043 37247
rect 29745 37213 29779 37247
rect 30573 37213 30607 37247
rect 31033 37213 31067 37247
rect 32597 37213 32631 37247
rect 33425 37213 33459 37247
rect 33609 37213 33643 37247
rect 34897 37213 34931 37247
rect 34989 37213 35023 37247
rect 36185 37213 36219 37247
rect 36369 37213 36403 37247
rect 36645 37213 36679 37247
rect 38301 37213 38335 37247
rect 39129 37213 39163 37247
rect 40049 37213 40083 37247
rect 40233 37213 40267 37247
rect 40325 37213 40359 37247
rect 40509 37213 40543 37247
rect 41521 37213 41555 37247
rect 41797 37213 41831 37247
rect 42257 37213 42291 37247
rect 42441 37213 42475 37247
rect 43453 37213 43487 37247
rect 46029 37213 46063 37247
rect 46305 37213 46339 37247
rect 46673 37213 46707 37247
rect 47501 37213 47535 37247
rect 47593 37213 47627 37247
rect 48237 37213 48271 37247
rect 48330 37213 48364 37247
rect 48702 37213 48736 37247
rect 49341 37213 49375 37247
rect 49525 37213 49559 37247
rect 50721 37213 50755 37247
rect 50905 37213 50939 37247
rect 53389 37213 53423 37247
rect 54125 37213 54159 37247
rect 54218 37213 54252 37247
rect 54493 37213 54527 37247
rect 54590 37213 54624 37247
rect 56057 37213 56091 37247
rect 28457 37145 28491 37179
rect 29193 37145 29227 37179
rect 32229 37145 32263 37179
rect 33793 37145 33827 37179
rect 35173 37145 35207 37179
rect 36829 37145 36863 37179
rect 41705 37145 41739 37179
rect 47777 37145 47811 37179
rect 48513 37145 48547 37179
rect 48605 37145 48639 37179
rect 53665 37145 53699 37179
rect 54401 37145 54435 37179
rect 28273 37077 28307 37111
rect 29837 37077 29871 37111
rect 37841 37077 37875 37111
rect 40693 37077 40727 37111
rect 42625 37077 42659 37111
rect 45293 37077 45327 37111
rect 48881 37077 48915 37111
rect 52285 37077 52319 37111
rect 52745 37077 52779 37111
rect 54769 37077 54803 37111
rect 57989 37077 58023 37111
rect 30021 36873 30055 36907
rect 34345 36873 34379 36907
rect 36001 36873 36035 36907
rect 38485 36873 38519 36907
rect 48237 36873 48271 36907
rect 50169 36873 50203 36907
rect 51457 36873 51491 36907
rect 56149 36873 56183 36907
rect 29009 36805 29043 36839
rect 32505 36805 32539 36839
rect 46673 36805 46707 36839
rect 50353 36805 50387 36839
rect 51917 36805 51951 36839
rect 52193 36805 52227 36839
rect 28917 36737 28951 36771
rect 29193 36737 29227 36771
rect 29929 36737 29963 36771
rect 30757 36737 30791 36771
rect 31125 36737 31159 36771
rect 31217 36737 31251 36771
rect 32689 36737 32723 36771
rect 33333 36737 33367 36771
rect 34437 36737 34471 36771
rect 35357 36737 35391 36771
rect 35541 36737 35575 36771
rect 35633 36737 35667 36771
rect 35725 36737 35759 36771
rect 36461 36737 36495 36771
rect 36645 36737 36679 36771
rect 38117 36737 38151 36771
rect 38945 36737 38979 36771
rect 39037 36737 39071 36771
rect 39129 36737 39163 36771
rect 39589 36737 39623 36771
rect 40233 36737 40267 36771
rect 41153 36737 41187 36771
rect 41429 36737 41463 36771
rect 41613 36737 41647 36771
rect 42901 36737 42935 36771
rect 44649 36737 44683 36771
rect 45293 36737 45327 36771
rect 45477 36737 45511 36771
rect 45569 36737 45603 36771
rect 46397 36737 46431 36771
rect 46765 36737 46799 36771
rect 49249 36737 49283 36771
rect 50077 36737 50111 36771
rect 52101 36737 52135 36771
rect 52290 36737 52324 36771
rect 53205 36737 53239 36771
rect 53297 36737 53331 36771
rect 53389 36737 53423 36771
rect 53573 36737 53607 36771
rect 54769 36737 54803 36771
rect 30665 36669 30699 36703
rect 34253 36669 34287 36703
rect 36553 36669 36587 36703
rect 38025 36669 38059 36703
rect 44465 36669 44499 36703
rect 46213 36669 46247 36703
rect 47777 36669 47811 36703
rect 49157 36669 49191 36703
rect 49617 36669 49651 36703
rect 52193 36669 52227 36703
rect 54861 36669 54895 36703
rect 29193 36601 29227 36635
rect 34805 36601 34839 36635
rect 40417 36601 40451 36635
rect 44833 36601 44867 36635
rect 48145 36601 48179 36635
rect 55689 36601 55723 36635
rect 32873 36533 32907 36567
rect 33517 36533 33551 36567
rect 39681 36533 39715 36567
rect 40969 36533 41003 36567
rect 43085 36533 43119 36567
rect 45293 36533 45327 36567
rect 50353 36533 50387 36567
rect 50813 36533 50847 36567
rect 52929 36533 52963 36567
rect 54125 36533 54159 36567
rect 55137 36533 55171 36567
rect 56701 36533 56735 36567
rect 57345 36533 57379 36567
rect 58081 36533 58115 36567
rect 29193 36329 29227 36363
rect 34897 36329 34931 36363
rect 41245 36329 41279 36363
rect 44649 36329 44683 36363
rect 29837 36261 29871 36295
rect 44373 36261 44407 36295
rect 47593 36261 47627 36295
rect 53113 36261 53147 36295
rect 30481 36193 30515 36227
rect 30941 36193 30975 36227
rect 32873 36193 32907 36227
rect 36093 36193 36127 36227
rect 41153 36193 41187 36227
rect 41981 36193 42015 36227
rect 42901 36193 42935 36227
rect 44189 36193 44223 36227
rect 44281 36193 44315 36227
rect 45753 36193 45787 36227
rect 48881 36193 48915 36227
rect 49709 36193 49743 36227
rect 52837 36193 52871 36227
rect 53941 36193 53975 36227
rect 28917 36125 28951 36159
rect 29745 36125 29779 36159
rect 30573 36125 30607 36159
rect 31033 36125 31067 36159
rect 32045 36125 32079 36159
rect 33517 36125 33551 36159
rect 33610 36125 33644 36159
rect 33982 36125 34016 36159
rect 35081 36125 35115 36159
rect 35357 36125 35391 36159
rect 36529 36125 36563 36159
rect 36645 36125 36679 36159
rect 37657 36125 37691 36159
rect 37750 36125 37784 36159
rect 37933 36125 37967 36159
rect 38122 36125 38156 36159
rect 38761 36125 38795 36159
rect 40049 36125 40083 36159
rect 40969 36125 41003 36159
rect 41889 36125 41923 36159
rect 42257 36125 42291 36159
rect 42441 36125 42475 36159
rect 43085 36125 43119 36159
rect 43177 36125 43211 36159
rect 43545 36125 43579 36159
rect 44005 36125 44039 36159
rect 44465 36125 44499 36159
rect 45569 36125 45603 36159
rect 46489 36125 46523 36159
rect 46765 36125 46799 36159
rect 47409 36125 47443 36159
rect 47593 36125 47627 36159
rect 48053 36125 48087 36159
rect 48237 36125 48271 36159
rect 49065 36125 49099 36159
rect 50353 36125 50387 36159
rect 50446 36125 50480 36159
rect 50629 36125 50663 36159
rect 50859 36125 50893 36159
rect 52745 36125 52779 36159
rect 54033 36125 54067 36159
rect 55873 36125 55907 36159
rect 56149 36125 56183 36159
rect 57437 36125 57471 36159
rect 57713 36125 57747 36159
rect 29193 36057 29227 36091
rect 33793 36057 33827 36091
rect 33885 36057 33919 36091
rect 37105 36057 37139 36091
rect 38025 36057 38059 36091
rect 41337 36057 41371 36091
rect 45661 36057 45695 36091
rect 46949 36057 46983 36091
rect 50721 36057 50755 36091
rect 29009 35989 29043 36023
rect 34161 35989 34195 36023
rect 35265 35989 35299 36023
rect 36185 35989 36219 36023
rect 36277 35989 36311 36023
rect 38301 35989 38335 36023
rect 39405 35989 39439 36023
rect 40233 35989 40267 36023
rect 45201 35989 45235 36023
rect 46581 35989 46615 36023
rect 48145 35989 48179 36023
rect 49249 35989 49283 36023
rect 50997 35989 51031 36023
rect 51641 35989 51675 36023
rect 54861 35989 54895 36023
rect 55505 35989 55539 36023
rect 57069 35989 57103 36023
rect 29101 35785 29135 35819
rect 32689 35785 32723 35819
rect 35449 35785 35483 35819
rect 35817 35785 35851 35819
rect 41521 35785 41555 35819
rect 42717 35785 42751 35819
rect 43085 35785 43119 35819
rect 44189 35785 44223 35819
rect 45017 35785 45051 35819
rect 45385 35785 45419 35819
rect 56333 35785 56367 35819
rect 30389 35717 30423 35751
rect 33609 35717 33643 35751
rect 38301 35717 38335 35751
rect 38485 35717 38519 35751
rect 49893 35717 49927 35751
rect 50629 35717 50663 35751
rect 54769 35717 54803 35751
rect 56793 35717 56827 35751
rect 57345 35717 57379 35751
rect 29009 35649 29043 35683
rect 29285 35649 29319 35683
rect 30113 35649 30147 35683
rect 31217 35649 31251 35683
rect 31401 35649 31435 35683
rect 31769 35649 31803 35683
rect 36277 35649 36311 35683
rect 37473 35649 37507 35683
rect 37565 35649 37599 35683
rect 37749 35649 37783 35683
rect 38577 35649 38611 35683
rect 39221 35649 39255 35683
rect 40233 35649 40267 35683
rect 41429 35649 41463 35683
rect 41613 35649 41647 35683
rect 42625 35649 42659 35683
rect 42901 35649 42935 35683
rect 44097 35649 44131 35683
rect 44925 35649 44959 35683
rect 45201 35649 45235 35683
rect 46029 35649 46063 35683
rect 46213 35649 46247 35683
rect 46305 35649 46339 35683
rect 46397 35649 46431 35683
rect 47225 35649 47259 35683
rect 47961 35649 47995 35683
rect 48789 35649 48823 35683
rect 49157 35649 49191 35683
rect 50353 35649 50387 35683
rect 50446 35649 50480 35683
rect 50721 35649 50755 35683
rect 50859 35649 50893 35683
rect 51641 35649 51675 35683
rect 53205 35649 53239 35683
rect 54493 35649 54527 35683
rect 54586 35649 54620 35683
rect 54861 35649 54895 35683
rect 54958 35649 54992 35683
rect 55965 35649 55999 35683
rect 32505 35581 32539 35615
rect 32873 35581 32907 35615
rect 34161 35581 34195 35615
rect 35265 35581 35299 35615
rect 35357 35581 35391 35615
rect 39129 35581 39163 35615
rect 40141 35581 40175 35615
rect 48053 35581 48087 35615
rect 48973 35581 49007 35615
rect 51549 35581 51583 35615
rect 53113 35581 53147 35615
rect 53941 35581 53975 35615
rect 55873 35581 55907 35615
rect 29285 35513 29319 35547
rect 37749 35513 37783 35547
rect 38301 35513 38335 35547
rect 39589 35513 39623 35547
rect 40601 35513 40635 35547
rect 48329 35513 48363 35547
rect 49157 35513 49191 35547
rect 50997 35513 51031 35547
rect 52009 35513 52043 35547
rect 55137 35513 55171 35547
rect 32321 35445 32355 35479
rect 36369 35445 36403 35479
rect 43637 35445 43671 35479
rect 46673 35445 46707 35479
rect 58081 35445 58115 35479
rect 29193 35241 29227 35275
rect 30665 35241 30699 35275
rect 33425 35241 33459 35275
rect 34897 35241 34931 35275
rect 35449 35241 35483 35275
rect 39313 35241 39347 35275
rect 47317 35241 47351 35275
rect 49709 35241 49743 35275
rect 52193 35241 52227 35275
rect 52745 35241 52779 35275
rect 53665 35241 53699 35275
rect 32781 35173 32815 35207
rect 34253 35173 34287 35207
rect 43729 35173 43763 35207
rect 49157 35173 49191 35207
rect 57897 35173 57931 35207
rect 28825 35105 28859 35139
rect 37197 35105 37231 35139
rect 38761 35105 38795 35139
rect 42717 35105 42751 35139
rect 50537 35105 50571 35139
rect 53573 35105 53607 35139
rect 54861 35105 54895 35139
rect 57437 35105 57471 35139
rect 29009 35037 29043 35071
rect 30481 35037 30515 35071
rect 30665 35037 30699 35071
rect 31309 35037 31343 35071
rect 32413 35037 32447 35071
rect 32781 35037 32815 35071
rect 32965 35037 32999 35071
rect 33701 35037 33735 35071
rect 35633 35037 35667 35071
rect 35909 35037 35943 35071
rect 37013 35037 37047 35071
rect 37289 35037 37323 35071
rect 37381 35037 37415 35071
rect 37565 35037 37599 35071
rect 38025 35037 38059 35071
rect 38209 35037 38243 35071
rect 38669 35037 38703 35071
rect 38853 35037 38887 35071
rect 40785 35037 40819 35071
rect 41705 35037 41739 35071
rect 41889 35037 41923 35071
rect 42073 35037 42107 35071
rect 42809 35037 42843 35071
rect 44005 35037 44039 35071
rect 46673 35037 46707 35071
rect 46766 35037 46800 35071
rect 46949 35037 46983 35071
rect 47179 35037 47213 35071
rect 48605 35037 48639 35071
rect 48881 35037 48915 35071
rect 49249 35037 49283 35071
rect 50813 35037 50847 35071
rect 53757 35037 53791 35071
rect 53849 35037 53883 35071
rect 55965 35037 55999 35071
rect 56149 35037 56183 35071
rect 56241 35037 56275 35071
rect 57161 35037 57195 35071
rect 57345 35037 57379 35071
rect 27813 34969 27847 35003
rect 31861 34969 31895 35003
rect 33425 34969 33459 35003
rect 33609 34969 33643 35003
rect 38117 34969 38151 35003
rect 40141 34969 40175 35003
rect 43729 34969 43763 35003
rect 47041 34969 47075 35003
rect 35817 34901 35851 34935
rect 36829 34901 36863 34935
rect 40969 34901 41003 34935
rect 42901 34901 42935 34935
rect 43269 34901 43303 34935
rect 43913 34901 43947 34935
rect 44465 34901 44499 34935
rect 45293 34901 45327 34935
rect 47869 34901 47903 34935
rect 51457 34901 51491 34935
rect 54309 34901 54343 34935
rect 55781 34901 55815 34935
rect 56977 34901 57011 34935
rect 27537 34697 27571 34731
rect 32505 34697 32539 34731
rect 42625 34697 42659 34731
rect 48789 34697 48823 34731
rect 58179 34697 58213 34731
rect 30113 34629 30147 34663
rect 35265 34629 35299 34663
rect 36829 34629 36863 34663
rect 40325 34629 40359 34663
rect 40877 34629 40911 34663
rect 44281 34629 44315 34663
rect 53113 34629 53147 34663
rect 58265 34629 58299 34663
rect 27353 34561 27387 34595
rect 31125 34561 31159 34595
rect 31309 34561 31343 34595
rect 31585 34561 31619 34595
rect 32321 34561 32355 34595
rect 33149 34561 33183 34595
rect 33793 34561 33827 34595
rect 34805 34561 34839 34595
rect 35449 34561 35483 34595
rect 35541 34561 35575 34595
rect 36277 34561 36311 34595
rect 37473 34561 37507 34595
rect 37565 34561 37599 34595
rect 38301 34561 38335 34595
rect 41705 34561 41739 34595
rect 43453 34561 43487 34595
rect 45017 34561 45051 34595
rect 46029 34561 46063 34595
rect 47041 34561 47075 34595
rect 47961 34561 47995 34595
rect 48513 34561 48547 34595
rect 48973 34561 49007 34595
rect 49341 34561 49375 34595
rect 50997 34561 51031 34595
rect 51733 34561 51767 34595
rect 52929 34561 52963 34595
rect 54033 34561 54067 34595
rect 55505 34561 55539 34595
rect 56333 34561 56367 34595
rect 56517 34561 56551 34595
rect 57161 34561 57195 34595
rect 58081 34561 58115 34595
rect 58357 34561 58391 34595
rect 28089 34493 28123 34527
rect 31769 34493 31803 34527
rect 33885 34493 33919 34527
rect 34713 34493 34747 34527
rect 37749 34493 37783 34527
rect 41061 34493 41095 34527
rect 43545 34493 43579 34527
rect 45109 34493 45143 34527
rect 45937 34493 45971 34527
rect 46857 34493 46891 34527
rect 47225 34493 47259 34527
rect 51641 34493 51675 34527
rect 53941 34493 53975 34527
rect 55597 34493 55631 34527
rect 55873 34493 55907 34527
rect 57069 34493 57103 34527
rect 33333 34425 33367 34459
rect 41521 34425 41555 34459
rect 45385 34425 45419 34459
rect 52101 34425 52135 34459
rect 28352 34357 28386 34391
rect 36185 34357 36219 34391
rect 37657 34357 37691 34391
rect 38564 34357 38598 34391
rect 43729 34357 43763 34391
rect 46305 34357 46339 34391
rect 47869 34357 47903 34391
rect 50445 34357 50479 34391
rect 53297 34357 53331 34391
rect 54401 34357 54435 34391
rect 56425 34357 56459 34391
rect 57437 34357 57471 34391
rect 28273 34153 28307 34187
rect 29101 34153 29135 34187
rect 29745 34153 29779 34187
rect 31235 34153 31269 34187
rect 33057 34153 33091 34187
rect 36645 34153 36679 34187
rect 39405 34153 39439 34187
rect 43269 34153 43303 34187
rect 48881 34153 48915 34187
rect 57713 34153 57747 34187
rect 44649 34085 44683 34119
rect 54217 34085 54251 34119
rect 31493 34017 31527 34051
rect 33425 34017 33459 34051
rect 34897 34017 34931 34051
rect 35173 34017 35207 34051
rect 37657 34017 37691 34051
rect 40325 34017 40359 34051
rect 42073 34017 42107 34051
rect 42349 34017 42383 34051
rect 44189 34017 44223 34051
rect 47225 34017 47259 34051
rect 47961 34017 47995 34051
rect 55781 34017 55815 34051
rect 29009 33949 29043 33983
rect 32045 33949 32079 33983
rect 32413 33949 32447 33983
rect 33241 33949 33275 33983
rect 33517 33949 33551 33983
rect 33609 33949 33643 33983
rect 33793 33949 33827 33983
rect 37473 33949 37507 33983
rect 39313 33949 39347 33983
rect 42809 33949 42843 33983
rect 43085 33949 43119 33983
rect 44281 33949 44315 33983
rect 45753 33949 45787 33983
rect 45845 33949 45879 33983
rect 46029 33949 46063 33983
rect 47133 33949 47167 33983
rect 48697 33949 48731 33983
rect 49433 33949 49467 33983
rect 49617 33949 49651 33983
rect 50997 33949 51031 33983
rect 51089 33949 51123 33983
rect 51917 33949 51951 33983
rect 52101 33949 52135 33983
rect 53205 33949 53239 33983
rect 53389 33949 53423 33983
rect 53481 33949 53515 33983
rect 54493 33949 54527 33983
rect 55965 33949 55999 33983
rect 56057 33949 56091 33983
rect 56241 33949 56275 33983
rect 56333 33949 56367 33983
rect 27629 33881 27663 33915
rect 28181 33881 28215 33915
rect 37565 33881 37599 33915
rect 38393 33881 38427 33915
rect 38761 33881 38795 33915
rect 45201 33881 45235 33915
rect 47041 33881 47075 33915
rect 48421 33881 48455 33915
rect 49525 33881 49559 33915
rect 54217 33881 54251 33915
rect 57621 33881 57655 33915
rect 37105 33813 37139 33847
rect 42901 33813 42935 33847
rect 46213 33813 46247 33847
rect 46673 33813 46707 33847
rect 48513 33813 48547 33847
rect 50813 33813 50847 33847
rect 51457 33813 51491 33847
rect 52009 33813 52043 33847
rect 53021 33813 53055 33847
rect 54401 33813 54435 33847
rect 56793 33813 56827 33847
rect 31493 33609 31527 33643
rect 33425 33609 33459 33643
rect 35357 33609 35391 33643
rect 41981 33609 42015 33643
rect 53573 33609 53607 33643
rect 54033 33609 54067 33643
rect 57437 33609 57471 33643
rect 32413 33541 32447 33575
rect 32781 33541 32815 33575
rect 39957 33541 39991 33575
rect 29745 33473 29779 33507
rect 33241 33473 33275 33507
rect 33425 33473 33459 33507
rect 34713 33473 34747 33507
rect 35173 33473 35207 33507
rect 36553 33473 36587 33507
rect 41429 33473 41463 33507
rect 42073 33473 42107 33507
rect 42993 33473 43027 33507
rect 43545 33473 43579 33507
rect 43637 33473 43671 33507
rect 44557 33473 44591 33507
rect 44649 33473 44683 33507
rect 44833 33473 44867 33507
rect 46029 33473 46063 33507
rect 48237 33473 48271 33507
rect 48513 33473 48547 33507
rect 48697 33473 48731 33507
rect 49985 33473 50019 33507
rect 50261 33473 50295 33507
rect 50445 33473 50479 33507
rect 51365 33473 51399 33507
rect 52193 33473 52227 33507
rect 52377 33473 52411 33507
rect 53205 33473 53239 33507
rect 53389 33473 53423 33507
rect 54217 33473 54251 33507
rect 54401 33473 54435 33507
rect 57069 33473 57103 33507
rect 57529 33473 57563 33507
rect 30021 33405 30055 33439
rect 36645 33405 36679 33439
rect 37933 33405 37967 33439
rect 38209 33405 38243 33439
rect 42717 33405 42751 33439
rect 48421 33405 48455 33439
rect 50169 33405 50203 33439
rect 50997 33405 51031 33439
rect 51273 33405 51307 33439
rect 53113 33405 53147 33439
rect 53297 33405 53331 33439
rect 54493 33405 54527 33439
rect 55505 33405 55539 33439
rect 58081 33405 58115 33439
rect 42809 33337 42843 33371
rect 45017 33337 45051 33371
rect 48605 33337 48639 33371
rect 50077 33337 50111 33371
rect 52285 33337 52319 33371
rect 56057 33337 56091 33371
rect 28733 33269 28767 33303
rect 29193 33269 29227 33303
rect 34529 33269 34563 33303
rect 36829 33269 36863 33303
rect 40417 33269 40451 33303
rect 41337 33269 41371 33303
rect 42901 33269 42935 33303
rect 46121 33269 46155 33303
rect 46949 33269 46983 33303
rect 48881 33269 48915 33303
rect 49801 33269 49835 33303
rect 54953 33269 54987 33303
rect 57253 33269 57287 33303
rect 29193 33065 29227 33099
rect 30573 33065 30607 33099
rect 33057 33065 33091 33099
rect 36553 33065 36587 33099
rect 39037 33065 39071 33099
rect 41889 33065 41923 33099
rect 48513 33065 48547 33099
rect 49801 33065 49835 33099
rect 50353 33065 50387 33099
rect 52285 33065 52319 33099
rect 54493 33065 54527 33099
rect 55505 33065 55539 33099
rect 56609 33065 56643 33099
rect 57529 33065 57563 33099
rect 58265 33065 58299 33099
rect 36093 32997 36127 33031
rect 37197 32997 37231 33031
rect 46673 32997 46707 33031
rect 31309 32929 31343 32963
rect 35449 32929 35483 32963
rect 40141 32929 40175 32963
rect 46213 32929 46247 32963
rect 47317 32929 47351 32963
rect 48973 32929 49007 32963
rect 50721 32929 50755 32963
rect 57161 32929 57195 32963
rect 58081 32929 58115 32963
rect 29929 32861 29963 32895
rect 30665 32861 30699 32895
rect 33793 32861 33827 32895
rect 35725 32861 35759 32895
rect 36737 32861 36771 32895
rect 37381 32861 37415 32895
rect 37473 32861 37507 32895
rect 37749 32861 37783 32895
rect 38945 32861 38979 32895
rect 42809 32861 42843 32895
rect 42993 32861 43027 32895
rect 43086 32839 43120 32873
rect 43211 32861 43245 32895
rect 44373 32861 44407 32895
rect 45201 32861 45235 32895
rect 46305 32861 46339 32895
rect 47409 32861 47443 32895
rect 48697 32861 48731 32895
rect 48789 32861 48823 32895
rect 49065 32861 49099 32895
rect 49617 32861 49651 32895
rect 49801 32861 49835 32895
rect 50537 32861 50571 32895
rect 51273 32861 51307 32895
rect 51733 32861 51767 32895
rect 52469 32861 52503 32895
rect 52561 32861 52595 32895
rect 52745 32861 52779 32895
rect 52837 32861 52871 32895
rect 53941 32861 53975 32895
rect 54033 32861 54067 32895
rect 54217 32861 54251 32895
rect 54309 32861 54343 32895
rect 55689 32861 55723 32895
rect 55781 32861 55815 32895
rect 55965 32861 55999 32895
rect 56057 32861 56091 32895
rect 57253 32861 57287 32895
rect 58357 32861 58391 32895
rect 31585 32793 31619 32827
rect 33701 32793 33735 32827
rect 35633 32793 35667 32827
rect 37565 32793 37599 32827
rect 40417 32793 40451 32827
rect 43453 32793 43487 32827
rect 29837 32725 29871 32759
rect 38301 32725 38335 32759
rect 44465 32725 44499 32759
rect 45293 32725 45327 32759
rect 47777 32725 47811 32759
rect 53297 32725 53331 32759
rect 58081 32725 58115 32759
rect 30941 32521 30975 32555
rect 32321 32521 32355 32555
rect 34713 32521 34747 32555
rect 35725 32521 35759 32555
rect 37565 32521 37599 32555
rect 38025 32521 38059 32555
rect 39129 32521 39163 32555
rect 40785 32521 40819 32555
rect 41797 32521 41831 32555
rect 43177 32521 43211 32555
rect 46029 32521 46063 32555
rect 46581 32521 46615 32555
rect 47225 32521 47259 32555
rect 49709 32521 49743 32555
rect 51549 32521 51583 32555
rect 52929 32521 52963 32555
rect 54217 32521 54251 32555
rect 56241 32521 56275 32555
rect 57253 32521 57287 32555
rect 28365 32453 28399 32487
rect 36553 32453 36587 32487
rect 38302 32453 38336 32487
rect 38393 32453 38427 32487
rect 39405 32453 39439 32487
rect 40509 32453 40543 32487
rect 41521 32453 41555 32487
rect 44005 32453 44039 32487
rect 51825 32453 51859 32487
rect 53573 32453 53607 32487
rect 54861 32453 54895 32487
rect 55689 32453 55723 32487
rect 30389 32385 30423 32419
rect 31033 32385 31067 32419
rect 31493 32385 31527 32419
rect 32505 32385 32539 32419
rect 35449 32385 35483 32419
rect 36461 32385 36495 32419
rect 36645 32385 36679 32419
rect 36783 32385 36817 32419
rect 38210 32385 38244 32419
rect 38511 32385 38545 32419
rect 38669 32385 38703 32419
rect 39313 32385 39347 32419
rect 39497 32385 39531 32419
rect 39615 32385 39649 32419
rect 40233 32385 40267 32419
rect 40417 32385 40451 32419
rect 40601 32385 40635 32419
rect 41245 32385 41279 32419
rect 41429 32385 41463 32419
rect 41613 32385 41647 32419
rect 42809 32385 42843 32419
rect 42993 32385 43027 32419
rect 43729 32385 43763 32419
rect 48053 32385 48087 32419
rect 49341 32385 49375 32419
rect 50721 32385 50755 32419
rect 50813 32385 50847 32419
rect 50905 32385 50939 32419
rect 51089 32385 51123 32419
rect 51687 32385 51721 32419
rect 51917 32385 51951 32419
rect 52045 32385 52079 32419
rect 52193 32385 52227 32419
rect 53113 32385 53147 32419
rect 53205 32385 53239 32419
rect 53481 32385 53515 32419
rect 54493 32385 54527 32419
rect 55597 32385 55631 32419
rect 55965 32385 55999 32419
rect 56057 32385 56091 32419
rect 56701 32385 56735 32419
rect 56793 32385 56827 32419
rect 56977 32385 57011 32419
rect 57069 32385 57103 32419
rect 30113 32317 30147 32351
rect 32965 32317 32999 32351
rect 33241 32317 33275 32351
rect 36277 32317 36311 32351
rect 36921 32317 36955 32351
rect 39773 32317 39807 32351
rect 45477 32317 45511 32351
rect 47777 32317 47811 32351
rect 49433 32317 49467 32351
rect 50445 32317 50479 32351
rect 54401 32317 54435 32351
rect 54769 32317 54803 32351
rect 47869 32249 47903 32283
rect 48237 32181 48271 32215
rect 58081 32181 58115 32215
rect 30389 31977 30423 32011
rect 31217 31977 31251 32011
rect 34161 31977 34195 32011
rect 35357 31977 35391 32011
rect 36553 31977 36587 32011
rect 38761 31977 38795 32011
rect 41153 31977 41187 32011
rect 41613 31977 41647 32011
rect 46949 31977 46983 32011
rect 48145 31977 48179 32011
rect 49433 31977 49467 32011
rect 50997 31977 51031 32011
rect 53757 31977 53791 32011
rect 56425 31977 56459 32011
rect 40049 31909 40083 31943
rect 43637 31909 43671 31943
rect 52469 31909 52503 31943
rect 57897 31909 57931 31943
rect 32965 31841 32999 31875
rect 33517 31841 33551 31875
rect 35817 31841 35851 31875
rect 36001 31841 36035 31875
rect 42165 31841 42199 31875
rect 45845 31841 45879 31875
rect 47961 31841 47995 31875
rect 48789 31841 48823 31875
rect 51549 31841 51583 31875
rect 52377 31841 52411 31875
rect 54769 31841 54803 31875
rect 55873 31841 55907 31875
rect 56241 31841 56275 31875
rect 29929 31773 29963 31807
rect 33609 31773 33643 31807
rect 34253 31773 34287 31807
rect 36737 31773 36771 31807
rect 36829 31773 36863 31807
rect 37197 31773 37231 31807
rect 37657 31773 37691 31807
rect 40233 31773 40267 31807
rect 40417 31773 40451 31807
rect 40601 31773 40635 31807
rect 42993 31773 43027 31807
rect 43177 31773 43211 31807
rect 44281 31773 44315 31807
rect 45937 31773 45971 31807
rect 48237 31773 48271 31807
rect 48697 31773 48731 31807
rect 48881 31773 48915 31807
rect 49341 31773 49375 31807
rect 50721 31773 50755 31807
rect 50997 31773 51031 31807
rect 51457 31773 51491 31807
rect 51641 31773 51675 31807
rect 52561 31773 52595 31807
rect 52653 31773 52687 31807
rect 53113 31773 53147 31807
rect 53261 31773 53295 31807
rect 53389 31773 53423 31807
rect 53578 31773 53612 31807
rect 55781 31773 55815 31807
rect 56149 31773 56183 31807
rect 56885 31773 56919 31807
rect 57069 31773 57103 31807
rect 57621 31773 57655 31807
rect 57713 31773 57747 31807
rect 32689 31705 32723 31739
rect 35725 31705 35759 31739
rect 36921 31705 36955 31739
rect 37059 31705 37093 31739
rect 40325 31705 40359 31739
rect 46029 31705 46063 31739
rect 50813 31705 50847 31739
rect 53481 31705 53515 31739
rect 54585 31705 54619 31739
rect 57897 31705 57931 31739
rect 29837 31637 29871 31671
rect 38301 31637 38335 31671
rect 39313 31637 39347 31671
rect 43085 31637 43119 31671
rect 44373 31637 44407 31671
rect 46397 31637 46431 31671
rect 47409 31637 47443 31671
rect 47961 31637 47995 31671
rect 28457 31433 28491 31467
rect 32413 31433 32447 31467
rect 35081 31433 35115 31467
rect 35909 31433 35943 31467
rect 38117 31433 38151 31467
rect 38669 31433 38703 31467
rect 46121 31433 46155 31467
rect 50721 31433 50755 31467
rect 50905 31433 50939 31467
rect 51733 31433 51767 31467
rect 55229 31433 55263 31467
rect 56425 31433 56459 31467
rect 29929 31365 29963 31399
rect 38837 31365 38871 31399
rect 39037 31365 39071 31399
rect 40233 31365 40267 31399
rect 40463 31365 40497 31399
rect 41199 31365 41233 31399
rect 41429 31365 41463 31399
rect 46029 31365 46063 31399
rect 54217 31365 54251 31399
rect 55873 31365 55907 31399
rect 30205 31297 30239 31331
rect 32505 31297 32539 31331
rect 33333 31297 33367 31331
rect 37473 31297 37507 31331
rect 40141 31297 40175 31331
rect 40325 31297 40359 31331
rect 41337 31297 41371 31331
rect 41521 31297 41555 31331
rect 43361 31297 43395 31331
rect 44097 31297 44131 31331
rect 45201 31297 45235 31331
rect 46949 31297 46983 31331
rect 47133 31297 47167 31331
rect 47777 31297 47811 31331
rect 49157 31297 49191 31331
rect 49341 31297 49375 31331
rect 50780 31297 50814 31331
rect 51549 31297 51583 31331
rect 51825 31297 51859 31331
rect 53205 31297 53239 31331
rect 54493 31297 54527 31331
rect 54585 31297 54619 31331
rect 56149 31297 56183 31331
rect 56885 31297 56919 31331
rect 56977 31297 57011 31331
rect 57161 31297 57195 31331
rect 57253 31297 57287 31331
rect 58357 31297 58391 31331
rect 33609 31229 33643 31263
rect 36001 31229 36035 31263
rect 36093 31229 36127 31263
rect 39957 31229 39991 31263
rect 40601 31229 40635 31263
rect 41061 31229 41095 31263
rect 44925 31229 44959 31263
rect 45937 31229 45971 31263
rect 47869 31229 47903 31263
rect 48973 31229 49007 31263
rect 50261 31229 50295 31263
rect 52285 31229 52319 31263
rect 54125 31229 54159 31263
rect 55781 31229 55815 31263
rect 56241 31229 56275 31263
rect 58081 31229 58115 31263
rect 42717 31161 42751 31195
rect 43177 31161 43211 31195
rect 46489 31161 46523 31195
rect 48145 31161 48179 31195
rect 50353 31161 50387 31195
rect 58265 31161 58299 31195
rect 35541 31093 35575 31127
rect 36737 31093 36771 31127
rect 37565 31093 37599 31127
rect 38853 31093 38887 31127
rect 41705 31093 41739 31127
rect 44005 31093 44039 31127
rect 46949 31093 46983 31127
rect 47777 31093 47811 31127
rect 51365 31093 51399 31127
rect 53021 31093 53055 31127
rect 54769 31093 54803 31127
rect 57437 31093 57471 31127
rect 58173 31093 58207 31127
rect 33701 30889 33735 30923
rect 39129 30889 39163 30923
rect 39313 30889 39347 30923
rect 43269 30889 43303 30923
rect 49433 30889 49467 30923
rect 53481 30889 53515 30923
rect 57529 30889 57563 30923
rect 38209 30821 38243 30855
rect 45937 30821 45971 30855
rect 29837 30753 29871 30787
rect 35449 30753 35483 30787
rect 40049 30753 40083 30787
rect 41521 30753 41555 30787
rect 47409 30753 47443 30787
rect 48789 30753 48823 30787
rect 48973 30753 49007 30787
rect 52469 30753 52503 30787
rect 54217 30753 54251 30787
rect 57253 30753 57287 30787
rect 1869 30685 1903 30719
rect 31861 30685 31895 30719
rect 33057 30685 33091 30719
rect 33885 30685 33919 30719
rect 36461 30685 36495 30719
rect 40233 30685 40267 30719
rect 40417 30685 40451 30719
rect 40693 30685 40727 30719
rect 43821 30685 43855 30719
rect 44005 30685 44039 30719
rect 45477 30685 45511 30719
rect 45753 30685 45787 30719
rect 46397 30685 46431 30719
rect 46489 30685 46523 30719
rect 46673 30685 46707 30719
rect 46765 30685 46799 30719
rect 47593 30685 47627 30719
rect 47685 30685 47719 30719
rect 47895 30685 47929 30719
rect 48053 30685 48087 30719
rect 49065 30685 49099 30719
rect 50721 30685 50755 30719
rect 50997 30685 51031 30719
rect 51181 30685 51215 30719
rect 52561 30685 52595 30719
rect 54309 30685 54343 30719
rect 55505 30685 55539 30719
rect 55597 30685 55631 30719
rect 55781 30685 55815 30719
rect 55873 30685 55907 30719
rect 57161 30685 57195 30719
rect 31585 30617 31619 30651
rect 35265 30617 35299 30651
rect 36737 30617 36771 30651
rect 38945 30617 38979 30651
rect 40325 30617 40359 30651
rect 40535 30617 40569 30651
rect 41797 30617 41831 30651
rect 47777 30617 47811 30651
rect 51365 30617 51399 30651
rect 52837 30617 52871 30651
rect 52929 30617 52963 30651
rect 54585 30617 54619 30651
rect 54677 30617 54711 30651
rect 57989 30617 58023 30651
rect 1685 30549 1719 30583
rect 2421 30549 2455 30583
rect 33241 30549 33275 30583
rect 34897 30549 34931 30583
rect 35357 30549 35391 30583
rect 39145 30549 39179 30583
rect 44189 30549 44223 30583
rect 45569 30549 45603 30583
rect 46949 30549 46983 30583
rect 52285 30549 52319 30583
rect 54033 30549 54067 30583
rect 56057 30549 56091 30583
rect 36369 30345 36403 30379
rect 47869 30345 47903 30379
rect 30849 30277 30883 30311
rect 33885 30277 33919 30311
rect 34897 30277 34931 30311
rect 37749 30277 37783 30311
rect 37959 30277 37993 30311
rect 40049 30277 40083 30311
rect 40279 30277 40313 30311
rect 41337 30277 41371 30311
rect 45201 30277 45235 30311
rect 48513 30277 48547 30311
rect 49709 30277 49743 30311
rect 50629 30277 50663 30311
rect 50997 30277 51031 30311
rect 54769 30277 54803 30311
rect 56333 30277 56367 30311
rect 58081 30277 58115 30311
rect 28825 30209 28859 30243
rect 29469 30209 29503 30243
rect 29929 30209 29963 30243
rect 30941 30209 30975 30243
rect 34161 30209 34195 30243
rect 34621 30209 34655 30243
rect 37657 30209 37691 30243
rect 37842 30209 37876 30243
rect 38117 30209 38151 30243
rect 38761 30209 38795 30243
rect 39957 30209 39991 30243
rect 40141 30209 40175 30243
rect 41199 30209 41233 30243
rect 41428 30209 41462 30243
rect 41520 30209 41554 30243
rect 43177 30209 43211 30243
rect 46305 30209 46339 30243
rect 46397 30209 46431 30243
rect 46581 30209 46615 30243
rect 46673 30209 46707 30243
rect 47133 30209 47167 30243
rect 47777 30209 47811 30243
rect 47961 30209 47995 30243
rect 48421 30209 48455 30243
rect 48605 30209 48639 30243
rect 49341 30209 49375 30243
rect 50537 30209 50571 30243
rect 50813 30209 50847 30243
rect 52009 30209 52043 30243
rect 52101 30209 52135 30243
rect 52285 30209 52319 30243
rect 52377 30209 52411 30243
rect 53205 30209 53239 30243
rect 53665 30209 53699 30243
rect 53757 30209 53791 30243
rect 53941 30209 53975 30243
rect 54033 30209 54067 30243
rect 56057 30209 56091 30243
rect 57161 30209 57195 30243
rect 37473 30141 37507 30175
rect 38945 30141 38979 30175
rect 40417 30141 40451 30175
rect 41061 30141 41095 30175
rect 41705 30141 41739 30175
rect 43453 30141 43487 30175
rect 49157 30141 49191 30175
rect 55229 30141 55263 30175
rect 55965 30141 55999 30175
rect 56425 30141 56459 30175
rect 57069 30141 57103 30175
rect 28641 30073 28675 30107
rect 30113 30073 30147 30107
rect 39773 30073 39807 30107
rect 49617 30073 49651 30107
rect 57529 30073 57563 30107
rect 31493 30005 31527 30039
rect 32413 30005 32447 30039
rect 38577 30005 38611 30039
rect 42625 30005 42659 30039
rect 46121 30005 46155 30039
rect 51825 30005 51859 30039
rect 53021 30005 53055 30039
rect 54217 30005 54251 30039
rect 55781 30005 55815 30039
rect 29837 29801 29871 29835
rect 32505 29801 32539 29835
rect 34989 29801 35023 29835
rect 36461 29801 36495 29835
rect 40785 29801 40819 29835
rect 44557 29801 44591 29835
rect 46397 29801 46431 29835
rect 46489 29801 46523 29835
rect 47225 29801 47259 29835
rect 49249 29801 49283 29835
rect 49433 29801 49467 29835
rect 37565 29733 37599 29767
rect 38669 29733 38703 29767
rect 45845 29733 45879 29767
rect 47869 29733 47903 29767
rect 31585 29665 31619 29699
rect 37105 29665 37139 29699
rect 37933 29665 37967 29699
rect 39037 29665 39071 29699
rect 41245 29665 41279 29699
rect 41429 29665 41463 29699
rect 41981 29665 42015 29699
rect 46581 29665 46615 29699
rect 47041 29665 47075 29699
rect 50997 29665 51031 29699
rect 51917 29665 51951 29699
rect 54125 29665 54159 29699
rect 54493 29665 54527 29699
rect 56977 29665 57011 29699
rect 57253 29665 57287 29699
rect 34897 29597 34931 29631
rect 36645 29597 36679 29631
rect 36829 29597 36863 29631
rect 37749 29597 37783 29631
rect 38853 29597 38887 29631
rect 40325 29597 40359 29631
rect 44005 29597 44039 29631
rect 44465 29597 44499 29631
rect 45201 29597 45235 29631
rect 45294 29597 45328 29631
rect 45666 29597 45700 29631
rect 46305 29597 46339 29631
rect 47317 29597 47351 29631
rect 48053 29597 48087 29631
rect 48145 29597 48179 29631
rect 50353 29597 50387 29631
rect 50537 29597 50571 29631
rect 52009 29597 52043 29631
rect 53113 29597 53147 29631
rect 53205 29597 53239 29631
rect 53389 29597 53423 29631
rect 53481 29597 53515 29631
rect 54217 29597 54251 29631
rect 55689 29597 55723 29631
rect 55781 29597 55815 29631
rect 56057 29597 56091 29631
rect 56885 29597 56919 29631
rect 58081 29597 58115 29631
rect 31309 29529 31343 29563
rect 33793 29529 33827 29563
rect 34345 29529 34379 29563
rect 36737 29529 36771 29563
rect 36947 29529 36981 29563
rect 40049 29529 40083 29563
rect 40233 29529 40267 29563
rect 42257 29529 42291 29563
rect 45477 29529 45511 29563
rect 45569 29529 45603 29563
rect 47869 29529 47903 29563
rect 49065 29529 49099 29563
rect 49265 29529 49299 29563
rect 54585 29529 54619 29563
rect 56149 29529 56183 29563
rect 35541 29461 35575 29495
rect 40325 29461 40359 29495
rect 41153 29461 41187 29495
rect 47041 29461 47075 29495
rect 50445 29461 50479 29495
rect 52377 29461 52411 29495
rect 52929 29461 52963 29495
rect 53941 29461 53975 29495
rect 55505 29461 55539 29495
rect 58265 29461 58299 29495
rect 30205 29257 30239 29291
rect 32689 29257 32723 29291
rect 36921 29257 36955 29291
rect 37841 29257 37875 29291
rect 39221 29257 39255 29291
rect 39865 29257 39899 29291
rect 41705 29257 41739 29291
rect 43453 29257 43487 29291
rect 58173 29257 58207 29291
rect 40141 29189 40175 29223
rect 40233 29189 40267 29223
rect 41429 29189 41463 29223
rect 48145 29189 48179 29223
rect 53849 29189 53883 29223
rect 56977 29189 57011 29223
rect 30113 29121 30147 29155
rect 30849 29121 30883 29155
rect 31769 29121 31803 29155
rect 32597 29121 32631 29155
rect 33425 29121 33459 29155
rect 35910 29111 35944 29145
rect 36012 29121 36046 29155
rect 36106 29121 36140 29155
rect 36231 29121 36265 29155
rect 38393 29121 38427 29155
rect 38853 29121 38887 29155
rect 39037 29121 39071 29155
rect 40049 29121 40083 29155
rect 40371 29121 40405 29155
rect 40509 29121 40543 29155
rect 41061 29121 41095 29155
rect 41219 29121 41253 29155
rect 41337 29121 41371 29155
rect 41521 29121 41555 29155
rect 42625 29121 42659 29155
rect 42809 29121 42843 29155
rect 42901 29121 42935 29155
rect 43545 29121 43579 29155
rect 45134 29121 45168 29155
rect 46673 29121 46707 29155
rect 46765 29121 46799 29155
rect 46949 29121 46983 29155
rect 47041 29121 47075 29155
rect 47784 29121 47818 29155
rect 47925 29121 47959 29155
rect 48053 29121 48087 29155
rect 48283 29121 48317 29155
rect 49433 29121 49467 29155
rect 49525 29121 49559 29155
rect 49709 29121 49743 29155
rect 49801 29121 49835 29155
rect 50721 29121 50755 29155
rect 51917 29121 51951 29155
rect 53021 29121 53055 29155
rect 53205 29121 53239 29155
rect 54033 29121 54067 29155
rect 55137 29121 55171 29155
rect 55229 29121 55263 29155
rect 55413 29121 55447 29155
rect 55505 29121 55539 29155
rect 55965 29121 55999 29155
rect 56057 29121 56091 29155
rect 56241 29121 56275 29155
rect 56333 29121 56367 29155
rect 57345 29121 57379 29155
rect 33701 29053 33735 29087
rect 35725 29053 35759 29087
rect 36369 29053 36403 29087
rect 38117 29053 38151 29087
rect 44097 29053 44131 29087
rect 44281 29053 44315 29087
rect 45017 29053 45051 29087
rect 45293 29053 45327 29087
rect 45937 29053 45971 29087
rect 50813 29053 50847 29087
rect 51089 29053 51123 29087
rect 51825 29053 51859 29087
rect 35173 28985 35207 29019
rect 44741 28985 44775 29019
rect 31677 28917 31711 28951
rect 38301 28917 38335 28951
rect 42717 28917 42751 28951
rect 46489 28917 46523 28951
rect 48421 28917 48455 28951
rect 49249 28917 49283 28951
rect 51549 28917 51583 28951
rect 53113 28917 53147 28951
rect 53665 28917 53699 28951
rect 54953 28917 54987 28951
rect 56517 28917 56551 28951
rect 30849 28713 30883 28747
rect 34345 28713 34379 28747
rect 34989 28713 35023 28747
rect 36829 28713 36863 28747
rect 37197 28713 37231 28747
rect 40049 28713 40083 28747
rect 40417 28713 40451 28747
rect 45201 28713 45235 28747
rect 48237 28713 48271 28747
rect 50353 28713 50387 28747
rect 55597 28713 55631 28747
rect 56057 28713 56091 28747
rect 51641 28645 51675 28679
rect 54401 28645 54435 28679
rect 32597 28577 32631 28611
rect 35725 28577 35759 28611
rect 37105 28577 37139 28611
rect 38025 28577 38059 28611
rect 44005 28577 44039 28611
rect 49157 28577 49191 28611
rect 49341 28577 49375 28611
rect 54861 28577 54895 28611
rect 57805 28577 57839 28611
rect 57897 28577 57931 28611
rect 33057 28509 33091 28543
rect 35081 28509 35115 28543
rect 35909 28509 35943 28543
rect 36001 28509 36035 28543
rect 36369 28509 36403 28543
rect 37381 28509 37415 28543
rect 38117 28509 38151 28543
rect 38209 28509 38243 28543
rect 38853 28509 38887 28543
rect 40049 28509 40083 28543
rect 40141 28509 40175 28543
rect 41245 28509 41279 28543
rect 41547 28509 41581 28543
rect 41705 28509 41739 28543
rect 42349 28509 42383 28543
rect 43269 28509 43303 28543
rect 44189 28509 44223 28543
rect 45339 28509 45373 28543
rect 45569 28509 45603 28543
rect 45697 28509 45731 28543
rect 45845 28509 45879 28543
rect 46305 28509 46339 28543
rect 46397 28509 46431 28543
rect 46581 28509 46615 28543
rect 47501 28509 47535 28543
rect 47593 28509 47627 28543
rect 48237 28509 48271 28543
rect 48421 28509 48455 28543
rect 49065 28509 49099 28543
rect 49433 28509 49467 28543
rect 50353 28509 50387 28543
rect 50537 28509 50571 28543
rect 50997 28509 51031 28543
rect 51181 28509 51215 28543
rect 52285 28509 52319 28543
rect 53389 28509 53423 28543
rect 53481 28509 53515 28543
rect 53691 28509 53725 28543
rect 53849 28509 53883 28543
rect 54769 28509 54803 28543
rect 57713 28509 57747 28543
rect 32321 28441 32355 28475
rect 36093 28441 36127 28475
rect 36231 28441 36265 28475
rect 38945 28441 38979 28475
rect 39129 28441 39163 28475
rect 41337 28441 41371 28475
rect 41429 28441 41463 28475
rect 44097 28441 44131 28475
rect 45477 28441 45511 28475
rect 52377 28441 52411 28475
rect 53573 28441 53607 28475
rect 33149 28373 33183 28407
rect 33701 28373 33735 28407
rect 38393 28373 38427 28407
rect 38853 28373 38887 28407
rect 41061 28373 41095 28407
rect 42165 28373 42199 28407
rect 43177 28373 43211 28407
rect 44557 28373 44591 28407
rect 46765 28373 46799 28407
rect 47777 28373 47811 28407
rect 49065 28373 49099 28407
rect 51089 28373 51123 28407
rect 53205 28373 53239 28407
rect 56609 28373 56643 28407
rect 57345 28373 57379 28407
rect 37565 28169 37599 28203
rect 38301 28169 38335 28203
rect 40141 28169 40175 28203
rect 41429 28169 41463 28203
rect 41797 28169 41831 28203
rect 45385 28169 45419 28203
rect 45753 28169 45787 28203
rect 52009 28169 52043 28203
rect 53665 28169 53699 28203
rect 54309 28169 54343 28203
rect 34345 28101 34379 28135
rect 34805 28101 34839 28135
rect 46857 28101 46891 28135
rect 53297 28101 53331 28135
rect 53481 28101 53515 28135
rect 54125 28101 54159 28135
rect 37749 28033 37783 28067
rect 38853 28033 38887 28067
rect 39773 28033 39807 28067
rect 42625 28033 42659 28067
rect 43913 28033 43947 28067
rect 44006 28033 44040 28067
rect 44189 28033 44223 28067
rect 44281 28033 44315 28067
rect 44419 28033 44453 28067
rect 46213 28033 46247 28067
rect 46397 28033 46431 28067
rect 46489 28033 46523 28067
rect 46627 28033 46661 28067
rect 47777 28033 47811 28067
rect 47961 28033 47995 28067
rect 48789 28033 48823 28067
rect 48973 28033 49007 28067
rect 49985 28033 50019 28067
rect 50077 28033 50111 28067
rect 51089 28033 51123 28067
rect 51365 28033 51399 28067
rect 51549 28033 51583 28067
rect 54401 28033 54435 28067
rect 55505 28033 55539 28067
rect 57161 28033 57195 28067
rect 58357 28033 58391 28067
rect 32321 27965 32355 27999
rect 32597 27965 32631 27999
rect 38577 27965 38611 27999
rect 39865 27965 39899 27999
rect 41245 27965 41279 27999
rect 41337 27965 41371 27999
rect 43269 27965 43303 27999
rect 45201 27965 45235 27999
rect 45293 27965 45327 27999
rect 50169 27965 50203 27999
rect 50261 27965 50295 27999
rect 55597 27965 55631 27999
rect 57253 27965 57287 27999
rect 58081 27965 58115 27999
rect 49157 27897 49191 27931
rect 54125 27897 54159 27931
rect 57529 27897 57563 27931
rect 58265 27897 58299 27931
rect 31769 27829 31803 27863
rect 36093 27829 36127 27863
rect 38761 27829 38795 27863
rect 39957 27829 39991 27863
rect 42717 27829 42751 27863
rect 44557 27829 44591 27863
rect 47869 27829 47903 27863
rect 48973 27829 49007 27863
rect 50445 27829 50479 27863
rect 50905 27829 50939 27863
rect 55873 27829 55907 27863
rect 56333 27829 56367 27863
rect 58173 27829 58207 27863
rect 32597 27625 32631 27659
rect 37105 27625 37139 27659
rect 38577 27625 38611 27659
rect 40049 27625 40083 27659
rect 40969 27625 41003 27659
rect 41968 27625 42002 27659
rect 43453 27625 43487 27659
rect 46581 27625 46615 27659
rect 51181 27625 51215 27659
rect 52377 27625 52411 27659
rect 35265 27557 35299 27591
rect 37289 27557 37323 27591
rect 38761 27557 38795 27591
rect 39497 27557 39531 27591
rect 40417 27557 40451 27591
rect 47501 27557 47535 27591
rect 48697 27557 48731 27591
rect 50721 27557 50755 27591
rect 53021 27557 53055 27591
rect 35725 27489 35759 27523
rect 35909 27489 35943 27523
rect 41705 27489 41739 27523
rect 51917 27489 51951 27523
rect 53113 27489 53147 27523
rect 54125 27489 54159 27523
rect 57253 27489 57287 27523
rect 57437 27489 57471 27523
rect 57713 27489 57747 27523
rect 32781 27421 32815 27455
rect 33793 27421 33827 27455
rect 35633 27421 35667 27455
rect 36737 27421 36771 27455
rect 37105 27421 37139 27455
rect 38209 27421 38243 27455
rect 39405 27421 39439 27455
rect 39497 27421 39531 27455
rect 40049 27421 40083 27455
rect 40233 27421 40267 27455
rect 41153 27421 41187 27455
rect 44097 27421 44131 27455
rect 45385 27421 45419 27455
rect 45661 27421 45695 27455
rect 46121 27421 46155 27455
rect 46397 27421 46431 27455
rect 47685 27421 47719 27455
rect 47869 27421 47903 27455
rect 48329 27421 48363 27455
rect 49157 27421 49191 27455
rect 49433 27421 49467 27455
rect 50353 27421 50387 27455
rect 50537 27421 50571 27455
rect 51457 27421 51491 27455
rect 51641 27421 51675 27455
rect 51825 27421 51859 27455
rect 52653 27421 52687 27455
rect 52745 27421 52779 27455
rect 53941 27421 53975 27455
rect 54769 27421 54803 27455
rect 54953 27421 54987 27455
rect 55873 27421 55907 27455
rect 56425 27421 56459 27455
rect 57529 27421 57563 27455
rect 57621 27421 57655 27455
rect 34345 27353 34379 27387
rect 39221 27353 39255 27387
rect 44557 27353 44591 27387
rect 45569 27353 45603 27387
rect 46213 27353 46247 27387
rect 48513 27353 48547 27387
rect 49525 27353 49559 27387
rect 52837 27353 52871 27387
rect 55689 27353 55723 27387
rect 33609 27285 33643 27319
rect 38577 27285 38611 27319
rect 43913 27285 43947 27319
rect 45201 27285 45235 27319
rect 51549 27285 51583 27319
rect 53573 27285 53607 27319
rect 54033 27285 54067 27319
rect 54953 27285 54987 27319
rect 55505 27285 55539 27319
rect 58265 27285 58299 27319
rect 35633 27081 35667 27115
rect 37473 27081 37507 27115
rect 39037 27081 39071 27115
rect 39589 27081 39623 27115
rect 45569 27081 45603 27115
rect 47869 27081 47903 27115
rect 54309 27081 54343 27115
rect 54769 27081 54803 27115
rect 55965 27081 55999 27115
rect 33425 27013 33459 27047
rect 36829 27013 36863 27047
rect 37933 27013 37967 27047
rect 42809 27013 42843 27047
rect 43913 27013 43947 27047
rect 55045 27013 55079 27047
rect 55137 27013 55171 27047
rect 55781 27013 55815 27047
rect 56609 27013 56643 27047
rect 36001 26945 36035 26979
rect 36093 26945 36127 26979
rect 38485 26945 38519 26979
rect 39497 26945 39531 26979
rect 39681 26945 39715 26979
rect 40693 26945 40727 26979
rect 41153 26945 41187 26979
rect 43085 26945 43119 26979
rect 43637 26945 43671 26979
rect 44557 26945 44591 26979
rect 44649 26945 44683 26979
rect 44833 26945 44867 26979
rect 46213 26945 46247 26979
rect 46397 26945 46431 26979
rect 47041 26945 47075 26979
rect 47225 26945 47259 26979
rect 47777 26945 47811 26979
rect 47961 26945 47995 26979
rect 48789 26945 48823 26979
rect 48973 26945 49007 26979
rect 50077 26945 50111 26979
rect 50169 26945 50203 26979
rect 50353 26945 50387 26979
rect 50445 26945 50479 26979
rect 50537 26945 50571 26979
rect 51365 26945 51399 26979
rect 51457 26945 51491 26979
rect 51733 26945 51767 26979
rect 53389 26945 53423 26979
rect 54953 26945 54987 26979
rect 55321 26945 55355 26979
rect 56057 26945 56091 26979
rect 33149 26877 33183 26911
rect 35173 26877 35207 26911
rect 36277 26877 36311 26911
rect 38761 26877 38795 26911
rect 53297 26877 53331 26911
rect 37565 26809 37599 26843
rect 46489 26809 46523 26843
rect 50721 26809 50755 26843
rect 53757 26809 53791 26843
rect 55781 26809 55815 26843
rect 38577 26741 38611 26775
rect 45017 26741 45051 26775
rect 47133 26741 47167 26775
rect 49157 26741 49191 26775
rect 51181 26741 51215 26775
rect 51641 26741 51675 26775
rect 52193 26741 52227 26775
rect 57161 26741 57195 26775
rect 58081 26741 58115 26775
rect 31677 26537 31711 26571
rect 34253 26537 34287 26571
rect 36645 26537 36679 26571
rect 37933 26537 37967 26571
rect 40049 26537 40083 26571
rect 40233 26537 40267 26571
rect 41889 26537 41923 26571
rect 45293 26537 45327 26571
rect 47041 26537 47075 26571
rect 50445 26537 50479 26571
rect 52377 26537 52411 26571
rect 52929 26537 52963 26571
rect 53573 26537 53607 26571
rect 54309 26537 54343 26571
rect 54677 26537 54711 26571
rect 55597 26537 55631 26571
rect 56701 26537 56735 26571
rect 42441 26469 42475 26503
rect 47869 26469 47903 26503
rect 56057 26469 56091 26503
rect 34897 26401 34931 26435
rect 37565 26401 37599 26435
rect 39221 26401 39255 26435
rect 40325 26401 40359 26435
rect 41337 26401 41371 26435
rect 44189 26401 44223 26435
rect 46489 26401 46523 26435
rect 48053 26401 48087 26435
rect 54217 26401 54251 26435
rect 32965 26333 32999 26367
rect 34161 26333 34195 26367
rect 37657 26333 37691 26367
rect 37749 26333 37783 26367
rect 39497 26333 39531 26367
rect 40601 26333 40635 26367
rect 41429 26333 41463 26367
rect 45201 26333 45235 26367
rect 47041 26333 47075 26367
rect 47225 26333 47259 26367
rect 47777 26333 47811 26367
rect 48513 26333 48547 26367
rect 48697 26333 48731 26367
rect 49157 26333 49191 26367
rect 49341 26333 49375 26367
rect 49433 26333 49467 26367
rect 49525 26333 49559 26367
rect 50353 26333 50387 26367
rect 50537 26333 50571 26367
rect 50997 26333 51031 26367
rect 51264 26333 51298 26367
rect 54493 26333 54527 26367
rect 35173 26265 35207 26299
rect 43913 26265 43947 26299
rect 46305 26265 46339 26299
rect 48053 26265 48087 26299
rect 49801 26265 49835 26299
rect 57253 26265 57287 26299
rect 41521 26197 41555 26231
rect 45845 26197 45879 26231
rect 46213 26197 46247 26231
rect 48697 26197 48731 26231
rect 34529 25993 34563 26027
rect 35173 25993 35207 26027
rect 37473 25993 37507 26027
rect 39589 25993 39623 26027
rect 43637 25993 43671 26027
rect 46305 25993 46339 26027
rect 46949 25993 46983 26027
rect 49709 25993 49743 26027
rect 50445 25993 50479 26027
rect 52101 25993 52135 26027
rect 53665 25993 53699 26027
rect 54585 25993 54619 26027
rect 55689 25993 55723 26027
rect 56241 25993 56275 26027
rect 36185 25925 36219 25959
rect 40141 25925 40175 25959
rect 42901 25925 42935 25959
rect 48053 25925 48087 25959
rect 49065 25925 49099 25959
rect 49249 25925 49283 25959
rect 50905 25925 50939 25959
rect 55229 25925 55263 25959
rect 34989 25857 35023 25891
rect 37657 25857 37691 25891
rect 37933 25857 37967 25891
rect 38393 25857 38427 25891
rect 38577 25857 38611 25891
rect 39313 25857 39347 25891
rect 39681 25857 39715 25891
rect 41061 25857 41095 25891
rect 41981 25857 42015 25891
rect 42625 25857 42659 25891
rect 43729 25857 43763 25891
rect 44465 25857 44499 25891
rect 46121 25857 46155 25891
rect 47961 25857 47995 25891
rect 48145 25857 48179 25891
rect 48329 25857 48363 25891
rect 48421 25857 48455 25891
rect 49709 25857 49743 25891
rect 49893 25857 49927 25891
rect 36277 25789 36311 25823
rect 36461 25789 36495 25823
rect 37841 25789 37875 25823
rect 39221 25789 39255 25823
rect 45937 25789 45971 25823
rect 35817 25721 35851 25755
rect 37933 25653 37967 25687
rect 38485 25653 38519 25687
rect 44281 25653 44315 25687
rect 44925 25653 44959 25687
rect 47777 25653 47811 25687
rect 48881 25653 48915 25687
rect 51549 25653 51583 25687
rect 35541 25449 35575 25483
rect 37473 25449 37507 25483
rect 38025 25449 38059 25483
rect 39129 25449 39163 25483
rect 39313 25449 39347 25483
rect 40509 25449 40543 25483
rect 43453 25449 43487 25483
rect 44005 25449 44039 25483
rect 44557 25449 44591 25483
rect 48237 25449 48271 25483
rect 49065 25449 49099 25483
rect 54401 25449 54435 25483
rect 38393 25381 38427 25415
rect 42901 25381 42935 25415
rect 47501 25381 47535 25415
rect 52653 25381 52687 25415
rect 40601 25313 40635 25347
rect 41153 25313 41187 25347
rect 47133 25313 47167 25347
rect 49709 25313 49743 25347
rect 51273 25313 51307 25347
rect 34345 25245 34379 25279
rect 35449 25245 35483 25279
rect 36461 25245 36495 25279
rect 38209 25245 38243 25279
rect 38485 25245 38519 25279
rect 38945 25245 38979 25279
rect 39037 25245 39071 25279
rect 40693 25245 40727 25279
rect 45201 25245 45235 25279
rect 46305 25245 46339 25279
rect 46489 25245 46523 25279
rect 47041 25245 47075 25279
rect 47225 25245 47259 25279
rect 47317 25245 47351 25279
rect 48329 25245 48363 25279
rect 48881 25245 48915 25279
rect 49157 25245 49191 25279
rect 50629 25245 50663 25279
rect 50813 25245 50847 25279
rect 36277 25177 36311 25211
rect 36645 25177 36679 25211
rect 37197 25177 37231 25211
rect 41429 25177 41463 25211
rect 48973 25177 49007 25211
rect 51518 25177 51552 25211
rect 34897 25109 34931 25143
rect 40325 25109 40359 25143
rect 45293 25109 45327 25143
rect 46305 25109 46339 25143
rect 50721 25109 50755 25143
rect 36369 24905 36403 24939
rect 37749 24837 37783 24871
rect 38853 24837 38887 24871
rect 39849 24837 39883 24871
rect 40049 24837 40083 24871
rect 41797 24837 41831 24871
rect 45845 24837 45879 24871
rect 34621 24769 34655 24803
rect 37657 24769 37691 24803
rect 37841 24769 37875 24803
rect 37979 24769 38013 24803
rect 38945 24769 38979 24803
rect 39221 24769 39255 24803
rect 40693 24769 40727 24803
rect 40877 24769 40911 24803
rect 41521 24769 41555 24803
rect 42809 24769 42843 24803
rect 42901 24769 42935 24803
rect 46489 24769 46523 24803
rect 46673 24769 46707 24803
rect 47869 24769 47903 24803
rect 48789 24769 48823 24803
rect 51181 24769 51215 24803
rect 51273 24769 51307 24803
rect 51549 24769 51583 24803
rect 34897 24701 34931 24735
rect 37473 24701 37507 24735
rect 38117 24701 38151 24735
rect 41797 24701 41831 24735
rect 42625 24701 42659 24735
rect 43821 24701 43855 24735
rect 44097 24701 44131 24735
rect 50997 24701 51031 24735
rect 51457 24701 51491 24735
rect 39681 24633 39715 24667
rect 41061 24633 41095 24667
rect 46857 24633 46891 24667
rect 39865 24565 39899 24599
rect 41613 24565 41647 24599
rect 42717 24565 42751 24599
rect 46673 24565 46707 24599
rect 50261 24565 50295 24599
rect 35817 24361 35851 24395
rect 42809 24361 42843 24395
rect 43453 24361 43487 24395
rect 44097 24361 44131 24395
rect 46489 24361 46523 24395
rect 49157 24361 49191 24395
rect 50813 24361 50847 24395
rect 36645 24293 36679 24327
rect 40141 24293 40175 24327
rect 37197 24225 37231 24259
rect 38025 24225 38059 24259
rect 40785 24225 40819 24259
rect 46305 24225 46339 24259
rect 47685 24225 47719 24259
rect 50445 24225 50479 24259
rect 35265 24157 35299 24191
rect 35909 24157 35943 24191
rect 38209 24157 38243 24191
rect 38301 24157 38335 24191
rect 39037 24157 39071 24191
rect 39405 24157 39439 24191
rect 39497 24157 39531 24191
rect 40049 24157 40083 24191
rect 40877 24157 40911 24191
rect 41521 24157 41555 24191
rect 41613 24157 41647 24191
rect 42717 24157 42751 24191
rect 43545 24157 43579 24191
rect 45201 24157 45235 24191
rect 46581 24157 46615 24191
rect 47409 24157 47443 24191
rect 50537 24157 50571 24191
rect 51365 24157 51399 24191
rect 37013 24089 37047 24123
rect 39129 24089 39163 24123
rect 39221 24089 39255 24123
rect 44649 24089 44683 24123
rect 35081 24021 35115 24055
rect 37105 24021 37139 24055
rect 38853 24021 38887 24055
rect 45293 24021 45327 24055
rect 46305 24021 46339 24055
rect 49709 24021 49743 24055
rect 51457 24021 51491 24055
rect 34345 23817 34379 23851
rect 36553 23817 36587 23851
rect 37933 23817 37967 23851
rect 39773 23817 39807 23851
rect 40325 23817 40359 23851
rect 47133 23817 47167 23851
rect 49157 23817 49191 23851
rect 35081 23749 35115 23783
rect 38117 23749 38151 23783
rect 44281 23749 44315 23783
rect 46029 23749 46063 23783
rect 49801 23749 49835 23783
rect 34805 23681 34839 23715
rect 37841 23681 37875 23715
rect 39221 23681 39255 23715
rect 42073 23681 42107 23715
rect 42809 23681 42843 23715
rect 43453 23681 43487 23715
rect 46489 23681 46523 23715
rect 47777 23681 47811 23715
rect 48053 23681 48087 23715
rect 49249 23681 49283 23715
rect 51825 23681 51859 23715
rect 41797 23613 41831 23647
rect 44005 23613 44039 23647
rect 51549 23613 51583 23647
rect 42625 23545 42659 23579
rect 43361 23545 43395 23579
rect 38117 23477 38151 23511
rect 46673 23477 46707 23511
rect 37841 23273 37875 23307
rect 39129 23273 39163 23307
rect 47961 23273 47995 23307
rect 51825 23273 51859 23307
rect 36001 23205 36035 23239
rect 44649 23205 44683 23239
rect 49341 23205 49375 23239
rect 37289 23137 37323 23171
rect 40049 23137 40083 23171
rect 46213 23137 46247 23171
rect 48881 23137 48915 23171
rect 36093 23069 36127 23103
rect 37197 23069 37231 23103
rect 37381 23069 37415 23103
rect 38669 23069 38703 23103
rect 39129 23069 39163 23103
rect 39405 23069 39439 23103
rect 42993 23069 43027 23103
rect 43821 23069 43855 23103
rect 44465 23069 44499 23103
rect 45385 23069 45419 23103
rect 48973 23069 49007 23103
rect 50353 23069 50387 23103
rect 40325 23001 40359 23035
rect 42073 23001 42107 23035
rect 42717 23001 42751 23035
rect 46489 23001 46523 23035
rect 38485 22933 38519 22967
rect 39313 22933 39347 22967
rect 43913 22933 43947 22967
rect 45201 22933 45235 22967
rect 36737 22729 36771 22763
rect 37565 22729 37599 22763
rect 39865 22729 39899 22763
rect 40785 22729 40819 22763
rect 41429 22729 41463 22763
rect 46673 22729 46707 22763
rect 49801 22729 49835 22763
rect 51089 22729 51123 22763
rect 44465 22661 44499 22695
rect 46213 22661 46247 22695
rect 36093 22593 36127 22627
rect 36921 22593 36955 22627
rect 37657 22593 37691 22627
rect 38117 22593 38151 22627
rect 40693 22593 40727 22627
rect 44189 22593 44223 22627
rect 46857 22593 46891 22627
rect 48053 22593 48087 22627
rect 50813 22593 50847 22627
rect 38393 22525 38427 22559
rect 48329 22525 48363 22559
rect 36277 22389 36311 22423
rect 51733 22389 51767 22423
rect 36264 22185 36298 22219
rect 48513 22185 48547 22219
rect 35449 22049 35483 22083
rect 36001 22049 36035 22083
rect 38025 22049 38059 22083
rect 38577 22049 38611 22083
rect 47317 22049 47351 22083
rect 49249 22049 49283 22083
rect 38485 21981 38519 22015
rect 38669 21981 38703 22015
rect 39313 21981 39347 22015
rect 47225 21981 47259 22015
rect 47869 21981 47903 22015
rect 48697 21981 48731 22015
rect 49341 21981 49375 22015
rect 39129 21845 39163 21879
rect 48053 21845 48087 21879
rect 37565 21641 37599 21675
rect 38301 21641 38335 21675
rect 39221 21641 39255 21675
rect 47777 21641 47811 21675
rect 37657 21505 37691 21539
rect 38117 21505 38151 21539
rect 39129 21505 39163 21539
rect 47317 21097 47351 21131
rect 48605 20893 48639 20927
rect 1593 2805 1627 2839
rect 58357 2805 58391 2839
rect 1777 2601 1811 2635
rect 29929 2601 29963 2635
rect 58173 2601 58207 2635
rect 1593 2397 1627 2431
rect 29745 2397 29779 2431
rect 58265 2329 58299 2363
rect 29101 2261 29135 2295
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 4874 57690
rect 4926 57638 4938 57690
rect 4990 57638 5002 57690
rect 5054 57638 5066 57690
rect 5118 57638 5130 57690
rect 5182 57638 35594 57690
rect 35646 57638 35658 57690
rect 35710 57638 35722 57690
rect 35774 57638 35786 57690
rect 35838 57638 35850 57690
rect 35902 57638 58880 57690
rect 1104 57616 58880 57638
rect 1302 57400 1308 57452
rect 1360 57440 1366 57452
rect 1581 57443 1639 57449
rect 1581 57440 1593 57443
rect 1360 57412 1593 57440
rect 1360 57400 1366 57412
rect 1581 57409 1593 57412
rect 1627 57440 1639 57443
rect 2961 57443 3019 57449
rect 2961 57440 2973 57443
rect 1627 57412 2973 57440
rect 1627 57409 1639 57412
rect 1581 57403 1639 57409
rect 2961 57409 2973 57412
rect 3007 57409 3019 57443
rect 2961 57403 3019 57409
rect 1765 57239 1823 57245
rect 1765 57205 1777 57239
rect 1811 57236 1823 57239
rect 1946 57236 1952 57248
rect 1811 57208 1952 57236
rect 1811 57205 1823 57208
rect 1765 57199 1823 57205
rect 1946 57196 1952 57208
rect 2004 57196 2010 57248
rect 2038 57196 2044 57248
rect 2096 57236 2102 57248
rect 2409 57239 2467 57245
rect 2409 57236 2421 57239
rect 2096 57208 2421 57236
rect 2096 57196 2102 57208
rect 2409 57205 2421 57208
rect 2455 57205 2467 57239
rect 2409 57199 2467 57205
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 2130 56896 2136 56908
rect 2091 56868 2136 56896
rect 2130 56856 2136 56868
rect 2188 56896 2194 56908
rect 2777 56899 2835 56905
rect 2777 56896 2789 56899
rect 2188 56868 2789 56896
rect 2188 56856 2194 56868
rect 2777 56865 2789 56868
rect 2823 56865 2835 56899
rect 2777 56859 2835 56865
rect 1946 56828 1952 56840
rect 1907 56800 1952 56828
rect 1946 56788 1952 56800
rect 2004 56788 2010 56840
rect 58253 56831 58311 56837
rect 58253 56797 58265 56831
rect 58299 56828 58311 56831
rect 58342 56828 58348 56840
rect 58299 56800 58348 56828
rect 58299 56797 58311 56800
rect 58253 56791 58311 56797
rect 58342 56788 58348 56800
rect 58400 56828 58406 56840
rect 59906 56828 59912 56840
rect 58400 56800 59912 56828
rect 58400 56788 58406 56800
rect 59906 56788 59912 56800
rect 59964 56788 59970 56840
rect 1578 56692 1584 56704
rect 1539 56664 1584 56692
rect 1578 56652 1584 56664
rect 1636 56652 1642 56704
rect 2038 56652 2044 56704
rect 2096 56692 2102 56704
rect 58161 56695 58219 56701
rect 2096 56664 2141 56692
rect 2096 56652 2102 56664
rect 58161 56661 58173 56695
rect 58207 56692 58219 56695
rect 58618 56692 58624 56704
rect 58207 56664 58624 56692
rect 58207 56661 58219 56664
rect 58161 56655 58219 56661
rect 58618 56652 58624 56664
rect 58676 56652 58682 56704
rect 1104 56602 58880 56624
rect 1104 56550 4874 56602
rect 4926 56550 4938 56602
rect 4990 56550 5002 56602
rect 5054 56550 5066 56602
rect 5118 56550 5130 56602
rect 5182 56550 35594 56602
rect 35646 56550 35658 56602
rect 35710 56550 35722 56602
rect 35774 56550 35786 56602
rect 35838 56550 35850 56602
rect 35902 56550 58880 56602
rect 1104 56528 58880 56550
rect 30374 56448 30380 56500
rect 30432 56488 30438 56500
rect 30926 56488 30932 56500
rect 30432 56460 30932 56488
rect 30432 56448 30438 56460
rect 30926 56448 30932 56460
rect 30984 56448 30990 56500
rect 58342 56488 58348 56500
rect 58303 56460 58348 56488
rect 58342 56448 58348 56460
rect 58400 56448 58406 56500
rect 1578 56380 1584 56432
rect 1636 56420 1642 56432
rect 1673 56423 1731 56429
rect 1673 56420 1685 56423
rect 1636 56392 1685 56420
rect 1636 56380 1642 56392
rect 1673 56389 1685 56392
rect 1719 56389 1731 56423
rect 1673 56383 1731 56389
rect 1949 56151 2007 56157
rect 1949 56117 1961 56151
rect 1995 56148 2007 56151
rect 2038 56148 2044 56160
rect 1995 56120 2044 56148
rect 1995 56117 2007 56120
rect 1949 56111 2007 56117
rect 2038 56108 2044 56120
rect 2096 56148 2102 56160
rect 30374 56148 30380 56160
rect 2096 56120 30380 56148
rect 2096 56108 2102 56120
rect 30374 56108 30380 56120
rect 30432 56108 30438 56160
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 1104 55514 58880 55536
rect 1104 55462 4874 55514
rect 4926 55462 4938 55514
rect 4990 55462 5002 55514
rect 5054 55462 5066 55514
rect 5118 55462 5130 55514
rect 5182 55462 35594 55514
rect 35646 55462 35658 55514
rect 35710 55462 35722 55514
rect 35774 55462 35786 55514
rect 35838 55462 35850 55514
rect 35902 55462 58880 55514
rect 1104 55440 58880 55462
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 1104 54426 58880 54448
rect 1104 54374 4874 54426
rect 4926 54374 4938 54426
rect 4990 54374 5002 54426
rect 5054 54374 5066 54426
rect 5118 54374 5130 54426
rect 5182 54374 35594 54426
rect 35646 54374 35658 54426
rect 35710 54374 35722 54426
rect 35774 54374 35786 54426
rect 35838 54374 35850 54426
rect 35902 54374 58880 54426
rect 1104 54352 58880 54374
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 1104 53338 58880 53360
rect 1104 53286 4874 53338
rect 4926 53286 4938 53338
rect 4990 53286 5002 53338
rect 5054 53286 5066 53338
rect 5118 53286 5130 53338
rect 5182 53286 35594 53338
rect 35646 53286 35658 53338
rect 35710 53286 35722 53338
rect 35774 53286 35786 53338
rect 35838 53286 35850 53338
rect 35902 53286 58880 53338
rect 1104 53264 58880 53286
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 1104 52250 58880 52272
rect 1104 52198 4874 52250
rect 4926 52198 4938 52250
rect 4990 52198 5002 52250
rect 5054 52198 5066 52250
rect 5118 52198 5130 52250
rect 5182 52198 35594 52250
rect 35646 52198 35658 52250
rect 35710 52198 35722 52250
rect 35774 52198 35786 52250
rect 35838 52198 35850 52250
rect 35902 52198 58880 52250
rect 1104 52176 58880 52198
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 1104 51162 58880 51184
rect 1104 51110 4874 51162
rect 4926 51110 4938 51162
rect 4990 51110 5002 51162
rect 5054 51110 5066 51162
rect 5118 51110 5130 51162
rect 5182 51110 35594 51162
rect 35646 51110 35658 51162
rect 35710 51110 35722 51162
rect 35774 51110 35786 51162
rect 35838 51110 35850 51162
rect 35902 51110 58880 51162
rect 1104 51088 58880 51110
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 4874 50074
rect 4926 50022 4938 50074
rect 4990 50022 5002 50074
rect 5054 50022 5066 50074
rect 5118 50022 5130 50074
rect 5182 50022 35594 50074
rect 35646 50022 35658 50074
rect 35710 50022 35722 50074
rect 35774 50022 35786 50074
rect 35838 50022 35850 50074
rect 35902 50022 58880 50074
rect 1104 50000 58880 50022
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1104 48986 58880 49008
rect 1104 48934 4874 48986
rect 4926 48934 4938 48986
rect 4990 48934 5002 48986
rect 5054 48934 5066 48986
rect 5118 48934 5130 48986
rect 5182 48934 35594 48986
rect 35646 48934 35658 48986
rect 35710 48934 35722 48986
rect 35774 48934 35786 48986
rect 35838 48934 35850 48986
rect 35902 48934 58880 48986
rect 1104 48912 58880 48934
rect 41785 48807 41843 48813
rect 36280 48776 38700 48804
rect 35342 48696 35348 48748
rect 35400 48736 35406 48748
rect 36173 48739 36231 48745
rect 36173 48736 36185 48739
rect 35400 48708 36185 48736
rect 35400 48696 35406 48708
rect 36173 48705 36185 48708
rect 36219 48705 36231 48739
rect 36173 48699 36231 48705
rect 36280 48680 36308 48776
rect 37642 48736 37648 48748
rect 37603 48708 37648 48736
rect 37642 48696 37648 48708
rect 37700 48696 37706 48748
rect 38672 48745 38700 48776
rect 41785 48773 41797 48807
rect 41831 48804 41843 48807
rect 43346 48804 43352 48816
rect 41831 48776 43352 48804
rect 41831 48773 41843 48776
rect 41785 48767 41843 48773
rect 43346 48764 43352 48776
rect 43404 48764 43410 48816
rect 38657 48739 38715 48745
rect 38657 48705 38669 48739
rect 38703 48705 38715 48739
rect 38657 48699 38715 48705
rect 39669 48739 39727 48745
rect 39669 48705 39681 48739
rect 39715 48736 39727 48739
rect 40218 48736 40224 48748
rect 39715 48708 40224 48736
rect 39715 48705 39727 48708
rect 39669 48699 39727 48705
rect 40218 48696 40224 48708
rect 40276 48696 40282 48748
rect 40586 48696 40592 48748
rect 40644 48736 40650 48748
rect 40773 48739 40831 48745
rect 40773 48736 40785 48739
rect 40644 48708 40785 48736
rect 40644 48696 40650 48708
rect 40773 48705 40785 48708
rect 40819 48705 40831 48739
rect 40954 48736 40960 48748
rect 40915 48708 40960 48736
rect 40773 48699 40831 48705
rect 40954 48696 40960 48708
rect 41012 48696 41018 48748
rect 42794 48736 42800 48748
rect 42755 48708 42800 48736
rect 42794 48696 42800 48708
rect 42852 48696 42858 48748
rect 43993 48739 44051 48745
rect 43993 48705 44005 48739
rect 44039 48705 44051 48739
rect 43993 48699 44051 48705
rect 36262 48668 36268 48680
rect 36175 48640 36268 48668
rect 36262 48628 36268 48640
rect 36320 48628 36326 48680
rect 37550 48668 37556 48680
rect 37511 48640 37556 48668
rect 37550 48628 37556 48640
rect 37608 48628 37614 48680
rect 38746 48668 38752 48680
rect 38707 48640 38752 48668
rect 38746 48628 38752 48640
rect 38804 48628 38810 48680
rect 39577 48671 39635 48677
rect 39577 48668 39589 48671
rect 39040 48640 39589 48668
rect 35345 48603 35403 48609
rect 35345 48600 35357 48603
rect 34256 48572 35357 48600
rect 34256 48544 34284 48572
rect 35345 48569 35357 48572
rect 35391 48569 35403 48603
rect 35345 48563 35403 48569
rect 36541 48603 36599 48609
rect 36541 48569 36553 48603
rect 36587 48600 36599 48603
rect 38470 48600 38476 48612
rect 36587 48572 38476 48600
rect 36587 48569 36599 48572
rect 36541 48563 36599 48569
rect 38470 48560 38476 48572
rect 38528 48560 38534 48612
rect 39040 48609 39068 48640
rect 39577 48637 39589 48640
rect 39623 48637 39635 48671
rect 39577 48631 39635 48637
rect 42889 48671 42947 48677
rect 42889 48637 42901 48671
rect 42935 48668 42947 48671
rect 44008 48668 44036 48699
rect 42935 48640 44036 48668
rect 44085 48671 44143 48677
rect 42935 48637 42947 48640
rect 42889 48631 42947 48637
rect 44085 48637 44097 48671
rect 44131 48637 44143 48671
rect 44085 48631 44143 48637
rect 39025 48603 39083 48609
rect 39025 48569 39037 48603
rect 39071 48569 39083 48603
rect 39025 48563 39083 48569
rect 40037 48603 40095 48609
rect 40037 48569 40049 48603
rect 40083 48600 40095 48603
rect 42904 48600 42932 48631
rect 40083 48572 42932 48600
rect 40083 48569 40095 48572
rect 40037 48563 40095 48569
rect 43346 48560 43352 48612
rect 43404 48600 43410 48612
rect 44100 48600 44128 48631
rect 43404 48572 44128 48600
rect 43404 48560 43410 48572
rect 33134 48492 33140 48544
rect 33192 48532 33198 48544
rect 33689 48535 33747 48541
rect 33689 48532 33701 48535
rect 33192 48504 33701 48532
rect 33192 48492 33198 48504
rect 33689 48501 33701 48504
rect 33735 48501 33747 48535
rect 34238 48532 34244 48544
rect 34199 48504 34244 48532
rect 33689 48495 33747 48501
rect 34238 48492 34244 48504
rect 34296 48492 34302 48544
rect 34790 48532 34796 48544
rect 34751 48504 34796 48532
rect 34790 48492 34796 48504
rect 34848 48492 34854 48544
rect 37921 48535 37979 48541
rect 37921 48501 37933 48535
rect 37967 48532 37979 48535
rect 38746 48532 38752 48544
rect 37967 48504 38752 48532
rect 37967 48501 37979 48504
rect 37921 48495 37979 48501
rect 38746 48492 38752 48504
rect 38804 48492 38810 48544
rect 43165 48535 43223 48541
rect 43165 48501 43177 48535
rect 43211 48532 43223 48535
rect 44266 48532 44272 48544
rect 43211 48504 44272 48532
rect 43211 48501 43223 48504
rect 43165 48495 43223 48501
rect 44266 48492 44272 48504
rect 44324 48492 44330 48544
rect 44358 48492 44364 48544
rect 44416 48532 44422 48544
rect 44416 48504 44461 48532
rect 44416 48492 44422 48504
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 35437 48263 35495 48269
rect 35437 48229 35449 48263
rect 35483 48260 35495 48263
rect 36262 48260 36268 48272
rect 35483 48232 36268 48260
rect 35483 48229 35495 48232
rect 35437 48223 35495 48229
rect 36262 48220 36268 48232
rect 36320 48220 36326 48272
rect 36449 48263 36507 48269
rect 36449 48229 36461 48263
rect 36495 48260 36507 48263
rect 37550 48260 37556 48272
rect 36495 48232 37556 48260
rect 36495 48229 36507 48232
rect 36449 48223 36507 48229
rect 37550 48220 37556 48232
rect 37608 48220 37614 48272
rect 38470 48220 38476 48272
rect 38528 48260 38534 48272
rect 40586 48260 40592 48272
rect 38528 48232 40264 48260
rect 40547 48232 40592 48260
rect 38528 48220 38534 48232
rect 33873 48195 33931 48201
rect 33873 48161 33885 48195
rect 33919 48161 33931 48195
rect 33873 48155 33931 48161
rect 34149 48195 34207 48201
rect 34149 48161 34161 48195
rect 34195 48192 34207 48195
rect 34977 48195 35035 48201
rect 34977 48192 34989 48195
rect 34195 48164 34989 48192
rect 34195 48161 34207 48164
rect 34149 48155 34207 48161
rect 34977 48161 34989 48164
rect 35023 48161 35035 48195
rect 35986 48192 35992 48204
rect 35947 48164 35992 48192
rect 34977 48155 35035 48161
rect 32582 48084 32588 48136
rect 32640 48124 32646 48136
rect 33781 48127 33839 48133
rect 33781 48124 33793 48127
rect 32640 48096 33793 48124
rect 32640 48084 32646 48096
rect 33781 48093 33793 48096
rect 33827 48093 33839 48127
rect 33781 48087 33839 48093
rect 33888 48056 33916 48155
rect 35986 48152 35992 48164
rect 36044 48152 36050 48204
rect 40126 48192 40132 48204
rect 40087 48164 40132 48192
rect 40126 48152 40132 48164
rect 40184 48152 40190 48204
rect 40236 48192 40264 48232
rect 40586 48220 40592 48232
rect 40644 48220 40650 48272
rect 41601 48263 41659 48269
rect 41601 48229 41613 48263
rect 41647 48260 41659 48263
rect 42886 48260 42892 48272
rect 41647 48232 42892 48260
rect 41647 48229 41659 48232
rect 41601 48223 41659 48229
rect 42886 48220 42892 48232
rect 42944 48220 42950 48272
rect 41141 48195 41199 48201
rect 41141 48192 41153 48195
rect 40236 48164 41153 48192
rect 41141 48161 41153 48164
rect 41187 48161 41199 48195
rect 41141 48155 41199 48161
rect 35066 48124 35072 48136
rect 35027 48096 35072 48124
rect 35066 48084 35072 48096
rect 35124 48084 35130 48136
rect 36081 48127 36139 48133
rect 36081 48093 36093 48127
rect 36127 48093 36139 48127
rect 36081 48087 36139 48093
rect 34698 48056 34704 48068
rect 33888 48028 34704 48056
rect 34698 48016 34704 48028
rect 34756 48056 34762 48068
rect 36096 48056 36124 48087
rect 38746 48084 38752 48136
rect 38804 48124 38810 48136
rect 40221 48127 40279 48133
rect 40221 48124 40233 48127
rect 38804 48096 40233 48124
rect 38804 48084 38810 48096
rect 40221 48093 40233 48096
rect 40267 48093 40279 48127
rect 41230 48124 41236 48136
rect 41191 48096 41236 48124
rect 40221 48087 40279 48093
rect 41230 48084 41236 48096
rect 41288 48084 41294 48136
rect 34756 48028 36124 48056
rect 34756 48016 34762 48028
rect 36722 48016 36728 48068
rect 36780 48056 36786 48068
rect 37001 48059 37059 48065
rect 37001 48056 37013 48059
rect 36780 48028 37013 48056
rect 36780 48016 36786 48028
rect 37001 48025 37013 48028
rect 37047 48056 37059 48059
rect 37553 48059 37611 48065
rect 37553 48056 37565 48059
rect 37047 48028 37565 48056
rect 37047 48025 37059 48028
rect 37001 48019 37059 48025
rect 37553 48025 37565 48028
rect 37599 48056 37611 48059
rect 37599 48028 38654 48056
rect 37599 48025 37611 48028
rect 37553 48019 37611 48025
rect 33134 47988 33140 48000
rect 33095 47960 33140 47988
rect 33134 47948 33140 47960
rect 33192 47948 33198 48000
rect 38105 47991 38163 47997
rect 38105 47957 38117 47991
rect 38151 47988 38163 47991
rect 38286 47988 38292 48000
rect 38151 47960 38292 47988
rect 38151 47957 38163 47960
rect 38105 47951 38163 47957
rect 38286 47948 38292 47960
rect 38344 47948 38350 48000
rect 38626 47988 38654 48028
rect 41782 47988 41788 48000
rect 38626 47960 41788 47988
rect 41782 47948 41788 47960
rect 41840 47988 41846 48000
rect 42061 47991 42119 47997
rect 42061 47988 42073 47991
rect 41840 47960 42073 47988
rect 41840 47948 41846 47960
rect 42061 47957 42073 47960
rect 42107 47957 42119 47991
rect 42061 47951 42119 47957
rect 1104 47898 58880 47920
rect 1104 47846 4874 47898
rect 4926 47846 4938 47898
rect 4990 47846 5002 47898
rect 5054 47846 5066 47898
rect 5118 47846 5130 47898
rect 5182 47846 35594 47898
rect 35646 47846 35658 47898
rect 35710 47846 35722 47898
rect 35774 47846 35786 47898
rect 35838 47846 35850 47898
rect 35902 47846 58880 47898
rect 1104 47824 58880 47846
rect 35066 47744 35072 47796
rect 35124 47784 35130 47796
rect 35618 47784 35624 47796
rect 35124 47756 35624 47784
rect 35124 47744 35130 47756
rect 35618 47744 35624 47756
rect 35676 47744 35682 47796
rect 39301 47787 39359 47793
rect 39301 47753 39313 47787
rect 39347 47784 39359 47787
rect 40126 47784 40132 47796
rect 39347 47756 40132 47784
rect 39347 47753 39359 47756
rect 39301 47747 39359 47753
rect 40126 47744 40132 47756
rect 40184 47744 40190 47796
rect 41325 47787 41383 47793
rect 41325 47753 41337 47787
rect 41371 47753 41383 47787
rect 41325 47747 41383 47753
rect 33134 47676 33140 47728
rect 33192 47716 33198 47728
rect 34885 47719 34943 47725
rect 34885 47716 34897 47719
rect 33192 47688 34897 47716
rect 33192 47676 33198 47688
rect 34885 47685 34897 47688
rect 34931 47716 34943 47719
rect 36078 47716 36084 47728
rect 34931 47688 36084 47716
rect 34931 47685 34943 47688
rect 34885 47679 34943 47685
rect 36078 47676 36084 47688
rect 36136 47716 36142 47728
rect 36633 47719 36691 47725
rect 36633 47716 36645 47719
rect 36136 47688 36645 47716
rect 36136 47676 36142 47688
rect 36633 47685 36645 47688
rect 36679 47685 36691 47719
rect 36633 47679 36691 47685
rect 32490 47648 32496 47660
rect 32451 47620 32496 47648
rect 32490 47608 32496 47620
rect 32548 47608 32554 47660
rect 33505 47651 33563 47657
rect 33505 47617 33517 47651
rect 33551 47617 33563 47651
rect 33505 47611 33563 47617
rect 32582 47580 32588 47592
rect 32543 47552 32588 47580
rect 32582 47540 32588 47552
rect 32640 47540 32646 47592
rect 32861 47583 32919 47589
rect 32861 47549 32873 47583
rect 32907 47580 32919 47583
rect 33413 47583 33471 47589
rect 33413 47580 33425 47583
rect 32907 47552 33425 47580
rect 32907 47549 32919 47552
rect 32861 47543 32919 47549
rect 33413 47549 33425 47552
rect 33459 47549 33471 47583
rect 33413 47543 33471 47549
rect 31662 47472 31668 47524
rect 31720 47512 31726 47524
rect 33520 47512 33548 47611
rect 35526 47608 35532 47660
rect 35584 47648 35590 47660
rect 35805 47651 35863 47657
rect 35805 47648 35817 47651
rect 35584 47620 35817 47648
rect 35584 47608 35590 47620
rect 35805 47617 35817 47620
rect 35851 47617 35863 47651
rect 35805 47611 35863 47617
rect 35986 47608 35992 47660
rect 36044 47648 36050 47660
rect 37645 47651 37703 47657
rect 37645 47648 37657 47651
rect 36044 47620 37657 47648
rect 36044 47608 36050 47620
rect 37645 47617 37657 47620
rect 37691 47617 37703 47651
rect 38930 47648 38936 47660
rect 38891 47620 38936 47648
rect 37645 47611 37703 47617
rect 38930 47608 38936 47620
rect 38988 47608 38994 47660
rect 40957 47651 41015 47657
rect 40957 47617 40969 47651
rect 41003 47617 41015 47651
rect 41340 47648 41368 47747
rect 42518 47648 42524 47660
rect 41340 47620 42524 47648
rect 40957 47611 41015 47617
rect 35713 47583 35771 47589
rect 35713 47549 35725 47583
rect 35759 47549 35771 47583
rect 37734 47580 37740 47592
rect 37695 47552 37740 47580
rect 35713 47543 35771 47549
rect 31720 47484 33548 47512
rect 33873 47515 33931 47521
rect 31720 47472 31726 47484
rect 33873 47481 33885 47515
rect 33919 47512 33931 47515
rect 35342 47512 35348 47524
rect 33919 47484 35348 47512
rect 33919 47481 33931 47484
rect 33873 47475 33931 47481
rect 35342 47472 35348 47484
rect 35400 47512 35406 47524
rect 35728 47512 35756 47543
rect 37734 47540 37740 47552
rect 37792 47540 37798 47592
rect 38841 47583 38899 47589
rect 38841 47580 38853 47583
rect 38028 47552 38853 47580
rect 38028 47521 38056 47552
rect 38841 47549 38853 47552
rect 38887 47549 38899 47583
rect 38841 47543 38899 47549
rect 40865 47583 40923 47589
rect 40865 47549 40877 47583
rect 40911 47549 40923 47583
rect 40972 47580 41000 47611
rect 42518 47608 42524 47620
rect 42576 47648 42582 47660
rect 42797 47651 42855 47657
rect 42797 47648 42809 47651
rect 42576 47620 42809 47648
rect 42576 47608 42582 47620
rect 42797 47617 42809 47620
rect 42843 47617 42855 47651
rect 44266 47648 44272 47660
rect 44227 47620 44272 47648
rect 42797 47611 42855 47617
rect 44266 47608 44272 47620
rect 44324 47608 44330 47660
rect 44450 47648 44456 47660
rect 44411 47620 44456 47648
rect 44450 47608 44456 47620
rect 44508 47608 44514 47660
rect 46474 47648 46480 47660
rect 46435 47620 46480 47648
rect 46474 47608 46480 47620
rect 46532 47608 46538 47660
rect 41414 47580 41420 47592
rect 40972 47552 41420 47580
rect 40865 47543 40923 47549
rect 35400 47484 35756 47512
rect 36173 47515 36231 47521
rect 35400 47472 35406 47484
rect 36173 47481 36185 47515
rect 36219 47512 36231 47515
rect 38013 47515 38071 47521
rect 36219 47484 37964 47512
rect 36219 47481 36231 47484
rect 36173 47475 36231 47481
rect 34514 47404 34520 47456
rect 34572 47444 34578 47456
rect 34609 47447 34667 47453
rect 34609 47444 34621 47447
rect 34572 47416 34621 47444
rect 34572 47404 34578 47416
rect 34609 47413 34621 47416
rect 34655 47413 34667 47447
rect 37936 47444 37964 47484
rect 38013 47481 38025 47515
rect 38059 47481 38071 47515
rect 40880 47512 40908 47543
rect 41414 47540 41420 47552
rect 41472 47540 41478 47592
rect 42886 47580 42892 47592
rect 42847 47552 42892 47580
rect 42886 47540 42892 47552
rect 42944 47540 42950 47592
rect 45281 47583 45339 47589
rect 45281 47549 45293 47583
rect 45327 47580 45339 47583
rect 45830 47580 45836 47592
rect 45327 47552 45836 47580
rect 45327 47549 45339 47552
rect 45281 47543 45339 47549
rect 45830 47540 45836 47552
rect 45888 47540 45894 47592
rect 46382 47580 46388 47592
rect 46343 47552 46388 47580
rect 46382 47540 46388 47552
rect 46440 47540 46446 47592
rect 38013 47475 38071 47481
rect 38488 47484 40908 47512
rect 38488 47444 38516 47484
rect 37936 47416 38516 47444
rect 34609 47407 34667 47413
rect 39758 47404 39764 47456
rect 39816 47444 39822 47456
rect 39853 47447 39911 47453
rect 39853 47444 39865 47447
rect 39816 47416 39865 47444
rect 39816 47404 39822 47416
rect 39853 47413 39865 47416
rect 39899 47444 39911 47447
rect 41874 47444 41880 47456
rect 39899 47416 41880 47444
rect 39899 47413 39911 47416
rect 39853 47407 39911 47413
rect 41874 47404 41880 47416
rect 41932 47404 41938 47456
rect 43070 47444 43076 47456
rect 43031 47416 43076 47444
rect 43070 47404 43076 47416
rect 43128 47404 43134 47456
rect 46845 47447 46903 47453
rect 46845 47413 46857 47447
rect 46891 47444 46903 47447
rect 47854 47444 47860 47456
rect 46891 47416 47860 47444
rect 46891 47413 46903 47416
rect 46845 47407 46903 47413
rect 47854 47404 47860 47416
rect 47912 47404 47918 47456
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 36817 47243 36875 47249
rect 36817 47240 36829 47243
rect 34164 47212 36829 47240
rect 32214 47132 32220 47184
rect 32272 47172 32278 47184
rect 34164 47181 34192 47212
rect 36817 47209 36829 47212
rect 36863 47240 36875 47243
rect 38013 47243 38071 47249
rect 38013 47240 38025 47243
rect 36863 47212 38025 47240
rect 36863 47209 36875 47212
rect 36817 47203 36875 47209
rect 38013 47209 38025 47212
rect 38059 47240 38071 47243
rect 38102 47240 38108 47252
rect 38059 47212 38108 47240
rect 38059 47209 38071 47212
rect 38013 47203 38071 47209
rect 38102 47200 38108 47212
rect 38160 47200 38166 47252
rect 34149 47175 34207 47181
rect 34149 47172 34161 47175
rect 32272 47144 34161 47172
rect 32272 47132 32278 47144
rect 34149 47141 34161 47144
rect 34195 47141 34207 47175
rect 34149 47135 34207 47141
rect 34348 47144 36676 47172
rect 32033 47107 32091 47113
rect 32033 47073 32045 47107
rect 32079 47104 32091 47107
rect 32858 47104 32864 47116
rect 32079 47076 32864 47104
rect 32079 47073 32091 47076
rect 32033 47067 32091 47073
rect 32858 47064 32864 47076
rect 32916 47104 32922 47116
rect 34348 47113 34376 47144
rect 36648 47113 36676 47144
rect 38470 47132 38476 47184
rect 38528 47172 38534 47184
rect 39301 47175 39359 47181
rect 39301 47172 39313 47175
rect 38528 47144 39313 47172
rect 38528 47132 38534 47144
rect 39301 47141 39313 47144
rect 39347 47141 39359 47175
rect 39301 47135 39359 47141
rect 40034 47132 40040 47184
rect 40092 47172 40098 47184
rect 41322 47172 41328 47184
rect 40092 47144 41328 47172
rect 40092 47132 40098 47144
rect 41322 47132 41328 47144
rect 41380 47132 41386 47184
rect 42981 47175 43039 47181
rect 42981 47141 42993 47175
rect 43027 47172 43039 47175
rect 45002 47172 45008 47184
rect 43027 47144 45008 47172
rect 43027 47141 43039 47144
rect 42981 47135 43039 47141
rect 45002 47132 45008 47144
rect 45060 47132 45066 47184
rect 45741 47175 45799 47181
rect 45741 47141 45753 47175
rect 45787 47172 45799 47175
rect 46382 47172 46388 47184
rect 45787 47144 46388 47172
rect 45787 47141 45799 47144
rect 45741 47135 45799 47141
rect 46382 47132 46388 47144
rect 46440 47132 46446 47184
rect 46753 47175 46811 47181
rect 46753 47141 46765 47175
rect 46799 47172 46811 47175
rect 47394 47172 47400 47184
rect 46799 47144 47400 47172
rect 46799 47141 46811 47144
rect 46753 47135 46811 47141
rect 47394 47132 47400 47144
rect 47452 47132 47458 47184
rect 34333 47107 34391 47113
rect 34333 47104 34345 47107
rect 32916 47076 34345 47104
rect 32916 47064 32922 47076
rect 34333 47073 34345 47076
rect 34379 47073 34391 47107
rect 34333 47067 34391 47073
rect 36633 47107 36691 47113
rect 36633 47073 36645 47107
rect 36679 47104 36691 47107
rect 37829 47107 37887 47113
rect 37829 47104 37841 47107
rect 36679 47076 37841 47104
rect 36679 47073 36691 47076
rect 36633 47067 36691 47073
rect 37829 47073 37841 47076
rect 37875 47104 37887 47107
rect 37918 47104 37924 47116
rect 37875 47076 37924 47104
rect 37875 47073 37887 47076
rect 37829 47067 37887 47073
rect 37918 47064 37924 47076
rect 37976 47064 37982 47116
rect 38841 47107 38899 47113
rect 38841 47073 38853 47107
rect 38887 47104 38899 47107
rect 39850 47104 39856 47116
rect 38887 47076 39856 47104
rect 38887 47073 38899 47076
rect 38841 47067 38899 47073
rect 39850 47064 39856 47076
rect 39908 47104 39914 47116
rect 40313 47107 40371 47113
rect 40313 47104 40325 47107
rect 39908 47076 40325 47104
rect 39908 47064 39914 47076
rect 40313 47073 40325 47076
rect 40359 47104 40371 47107
rect 40773 47107 40831 47113
rect 40773 47104 40785 47107
rect 40359 47076 40785 47104
rect 40359 47073 40371 47076
rect 40313 47067 40371 47073
rect 40773 47073 40785 47076
rect 40819 47073 40831 47107
rect 42518 47104 42524 47116
rect 42479 47076 42524 47104
rect 40773 47067 40831 47073
rect 42518 47064 42524 47076
rect 42576 47064 42582 47116
rect 43070 47064 43076 47116
rect 43128 47104 43134 47116
rect 45281 47107 45339 47113
rect 45281 47104 45293 47107
rect 43128 47076 45293 47104
rect 43128 47064 43134 47076
rect 45281 47073 45293 47076
rect 45327 47073 45339 47107
rect 45281 47067 45339 47073
rect 45830 47064 45836 47116
rect 45888 47104 45894 47116
rect 46293 47107 46351 47113
rect 46293 47104 46305 47107
rect 45888 47076 46305 47104
rect 45888 47064 45894 47076
rect 46293 47073 46305 47076
rect 46339 47073 46351 47107
rect 46293 47067 46351 47073
rect 32214 47036 32220 47048
rect 32175 47008 32220 47036
rect 32214 46996 32220 47008
rect 32272 46996 32278 47048
rect 32309 47039 32367 47045
rect 32309 47005 32321 47039
rect 32355 47036 32367 47039
rect 32674 47036 32680 47048
rect 32355 47008 32680 47036
rect 32355 47005 32367 47008
rect 32309 46999 32367 47005
rect 32674 46996 32680 47008
rect 32732 46996 32738 47048
rect 34057 47039 34115 47045
rect 34057 47005 34069 47039
rect 34103 47005 34115 47039
rect 34057 46999 34115 47005
rect 34885 47039 34943 47045
rect 34885 47005 34897 47039
rect 34931 47005 34943 47039
rect 34885 46999 34943 47005
rect 34978 47039 35036 47045
rect 34978 47005 34990 47039
rect 35024 47005 35036 47039
rect 34978 46999 35036 47005
rect 32122 46928 32128 46980
rect 32180 46968 32186 46980
rect 32861 46971 32919 46977
rect 32861 46968 32873 46971
rect 32180 46940 32873 46968
rect 32180 46928 32186 46940
rect 32861 46937 32873 46940
rect 32907 46937 32919 46971
rect 32861 46931 32919 46937
rect 33413 46971 33471 46977
rect 33413 46937 33425 46971
rect 33459 46968 33471 46971
rect 34072 46968 34100 46999
rect 33459 46940 34100 46968
rect 34333 46971 34391 46977
rect 33459 46937 33471 46940
rect 33413 46931 33471 46937
rect 34333 46937 34345 46971
rect 34379 46968 34391 46971
rect 34900 46968 34928 46999
rect 34379 46940 34928 46968
rect 34379 46937 34391 46940
rect 34333 46931 34391 46937
rect 32033 46903 32091 46909
rect 32033 46869 32045 46903
rect 32079 46900 32091 46903
rect 32306 46900 32312 46912
rect 32079 46872 32312 46900
rect 32079 46869 32091 46872
rect 32033 46863 32091 46869
rect 32306 46860 32312 46872
rect 32364 46860 32370 46912
rect 32950 46860 32956 46912
rect 33008 46900 33014 46912
rect 33134 46900 33140 46912
rect 33008 46872 33140 46900
rect 33008 46860 33014 46872
rect 33134 46860 33140 46872
rect 33192 46900 33198 46912
rect 33428 46900 33456 46931
rect 33192 46872 33456 46900
rect 33192 46860 33198 46872
rect 34514 46860 34520 46912
rect 34572 46900 34578 46912
rect 34992 46900 35020 46999
rect 35342 46996 35348 47048
rect 35400 47045 35406 47048
rect 35400 47036 35408 47045
rect 36081 47039 36139 47045
rect 35400 47008 35445 47036
rect 35400 46999 35408 47008
rect 36081 47005 36093 47039
rect 36127 47036 36139 47039
rect 36170 47036 36176 47048
rect 36127 47008 36176 47036
rect 36127 47005 36139 47008
rect 36081 46999 36139 47005
rect 35400 46996 35406 46999
rect 36170 46996 36176 47008
rect 36228 46996 36234 47048
rect 36722 47036 36728 47048
rect 36556 47008 36728 47036
rect 35158 46968 35164 46980
rect 35119 46940 35164 46968
rect 35158 46928 35164 46940
rect 35216 46928 35222 46980
rect 35253 46971 35311 46977
rect 35253 46937 35265 46971
rect 35299 46968 35311 46971
rect 36556 46968 36584 47008
rect 36722 46996 36728 47008
rect 36780 46996 36786 47048
rect 36909 47039 36967 47045
rect 36909 47005 36921 47039
rect 36955 47036 36967 47039
rect 37550 47036 37556 47048
rect 36955 47008 37556 47036
rect 36955 47005 36967 47008
rect 36909 46999 36967 47005
rect 37550 46996 37556 47008
rect 37608 46996 37614 47048
rect 38105 47039 38163 47045
rect 38105 47005 38117 47039
rect 38151 47005 38163 47039
rect 38105 46999 38163 47005
rect 38565 47039 38623 47045
rect 38565 47005 38577 47039
rect 38611 47005 38623 47039
rect 38565 46999 38623 47005
rect 38657 47039 38715 47045
rect 38657 47005 38669 47039
rect 38703 47036 38715 47039
rect 39298 47036 39304 47048
rect 38703 47008 39304 47036
rect 38703 47005 38715 47008
rect 38657 46999 38715 47005
rect 35299 46940 36584 46968
rect 36633 46971 36691 46977
rect 35299 46937 35311 46940
rect 35253 46931 35311 46937
rect 36633 46937 36645 46971
rect 36679 46968 36691 46971
rect 37458 46968 37464 46980
rect 36679 46940 37464 46968
rect 36679 46937 36691 46940
rect 36633 46931 36691 46937
rect 37458 46928 37464 46940
rect 37516 46928 37522 46980
rect 38120 46968 38148 46999
rect 38580 46968 38608 46999
rect 39298 46996 39304 47008
rect 39356 46996 39362 47048
rect 40034 47036 40040 47048
rect 39995 47008 40040 47036
rect 40034 46996 40040 47008
rect 40092 46996 40098 47048
rect 40129 47039 40187 47045
rect 40129 47005 40141 47039
rect 40175 47036 40187 47039
rect 40957 47039 41015 47045
rect 40957 47036 40969 47039
rect 40175 47008 40969 47036
rect 40175 47005 40187 47008
rect 40129 46999 40187 47005
rect 40957 47005 40969 47008
rect 41003 47005 41015 47039
rect 40957 46999 41015 47005
rect 41049 47039 41107 47045
rect 41049 47005 41061 47039
rect 41095 47036 41107 47039
rect 42613 47039 42671 47045
rect 41095 47008 41414 47036
rect 41095 47005 41107 47008
rect 41049 46999 41107 47005
rect 38746 46968 38752 46980
rect 38120 46940 38752 46968
rect 38746 46928 38752 46940
rect 38804 46928 38810 46980
rect 39316 46968 39344 46996
rect 40144 46968 40172 46999
rect 39316 46940 40172 46968
rect 34572 46872 35020 46900
rect 35529 46903 35587 46909
rect 34572 46860 34578 46872
rect 35529 46869 35541 46903
rect 35575 46900 35587 46903
rect 35618 46900 35624 46912
rect 35575 46872 35624 46900
rect 35575 46869 35587 46872
rect 35529 46863 35587 46869
rect 35618 46860 35624 46872
rect 35676 46860 35682 46912
rect 37829 46903 37887 46909
rect 37829 46869 37841 46903
rect 37875 46900 37887 46903
rect 38562 46900 38568 46912
rect 37875 46872 38568 46900
rect 37875 46869 37887 46872
rect 37829 46863 37887 46869
rect 38562 46860 38568 46872
rect 38620 46860 38626 46912
rect 38841 46903 38899 46909
rect 38841 46869 38853 46903
rect 38887 46900 38899 46903
rect 39206 46900 39212 46912
rect 38887 46872 39212 46900
rect 38887 46869 38899 46872
rect 38841 46863 38899 46869
rect 39206 46860 39212 46872
rect 39264 46860 39270 46912
rect 40310 46900 40316 46912
rect 40271 46872 40316 46900
rect 40310 46860 40316 46872
rect 40368 46860 40374 46912
rect 40402 46860 40408 46912
rect 40460 46900 40466 46912
rect 40773 46903 40831 46909
rect 40773 46900 40785 46903
rect 40460 46872 40785 46900
rect 40460 46860 40466 46872
rect 40773 46869 40785 46872
rect 40819 46869 40831 46903
rect 41386 46900 41414 47008
rect 42613 47005 42625 47039
rect 42659 47036 42671 47039
rect 43254 47036 43260 47048
rect 42659 47008 43260 47036
rect 42659 47005 42671 47008
rect 42613 46999 42671 47005
rect 43254 46996 43260 47008
rect 43312 46996 43318 47048
rect 45370 47036 45376 47048
rect 45331 47008 45376 47036
rect 45370 46996 45376 47008
rect 45428 46996 45434 47048
rect 46400 47045 46428 47132
rect 46385 47039 46443 47045
rect 46385 47005 46397 47039
rect 46431 47005 46443 47039
rect 46385 46999 46443 47005
rect 41506 46900 41512 46912
rect 41386 46872 41512 46900
rect 40773 46863 40831 46869
rect 41506 46860 41512 46872
rect 41564 46860 41570 46912
rect 41601 46903 41659 46909
rect 41601 46869 41613 46903
rect 41647 46900 41659 46903
rect 42978 46900 42984 46912
rect 41647 46872 42984 46900
rect 41647 46869 41659 46872
rect 41601 46863 41659 46869
rect 42978 46860 42984 46872
rect 43036 46900 43042 46912
rect 43533 46903 43591 46909
rect 43533 46900 43545 46903
rect 43036 46872 43545 46900
rect 43036 46860 43042 46872
rect 43533 46869 43545 46872
rect 43579 46900 43591 46903
rect 43993 46903 44051 46909
rect 43993 46900 44005 46903
rect 43579 46872 44005 46900
rect 43579 46869 43591 46872
rect 43533 46863 43591 46869
rect 43993 46869 44005 46872
rect 44039 46869 44051 46903
rect 44634 46900 44640 46912
rect 44595 46872 44640 46900
rect 43993 46863 44051 46869
rect 44634 46860 44640 46872
rect 44692 46860 44698 46912
rect 1104 46810 58880 46832
rect 1104 46758 4874 46810
rect 4926 46758 4938 46810
rect 4990 46758 5002 46810
rect 5054 46758 5066 46810
rect 5118 46758 5130 46810
rect 5182 46758 35594 46810
rect 35646 46758 35658 46810
rect 35710 46758 35722 46810
rect 35774 46758 35786 46810
rect 35838 46758 35850 46810
rect 35902 46758 58880 46810
rect 1104 46736 58880 46758
rect 32582 46696 32588 46708
rect 32543 46668 32588 46696
rect 32582 46656 32588 46668
rect 32640 46656 32646 46708
rect 34698 46696 34704 46708
rect 34659 46668 34704 46696
rect 34698 46656 34704 46668
rect 34756 46656 34762 46708
rect 37642 46656 37648 46708
rect 37700 46696 37706 46708
rect 38105 46699 38163 46705
rect 38105 46696 38117 46699
rect 37700 46668 38117 46696
rect 37700 46656 37706 46668
rect 38105 46665 38117 46668
rect 38151 46665 38163 46699
rect 38105 46659 38163 46665
rect 38746 46656 38752 46708
rect 38804 46656 38810 46708
rect 38930 46656 38936 46708
rect 38988 46696 38994 46708
rect 39209 46699 39267 46705
rect 39209 46696 39221 46699
rect 38988 46668 39221 46696
rect 38988 46656 38994 46668
rect 39209 46665 39221 46668
rect 39255 46665 39267 46699
rect 39209 46659 39267 46665
rect 40218 46656 40224 46708
rect 40276 46696 40282 46708
rect 40313 46699 40371 46705
rect 40313 46696 40325 46699
rect 40276 46668 40325 46696
rect 40276 46656 40282 46668
rect 40313 46665 40325 46668
rect 40359 46665 40371 46699
rect 40313 46659 40371 46665
rect 40770 46656 40776 46708
rect 40828 46696 40834 46708
rect 40828 46668 41276 46696
rect 40828 46656 40834 46668
rect 31205 46631 31263 46637
rect 31205 46597 31217 46631
rect 31251 46628 31263 46631
rect 34238 46628 34244 46640
rect 31251 46600 34244 46628
rect 31251 46597 31263 46600
rect 31205 46591 31263 46597
rect 31754 46520 31760 46572
rect 31812 46560 31818 46572
rect 33244 46569 33272 46600
rect 34238 46588 34244 46600
rect 34296 46588 34302 46640
rect 35158 46588 35164 46640
rect 35216 46628 35222 46640
rect 38764 46628 38792 46656
rect 40037 46631 40095 46637
rect 40037 46628 40049 46631
rect 35216 46600 37780 46628
rect 38764 46600 40049 46628
rect 35216 46588 35222 46600
rect 32309 46563 32367 46569
rect 32309 46560 32321 46563
rect 31812 46532 32321 46560
rect 31812 46520 31818 46532
rect 32309 46529 32321 46532
rect 32355 46529 32367 46563
rect 32309 46523 32367 46529
rect 33229 46563 33287 46569
rect 33229 46529 33241 46563
rect 33275 46529 33287 46563
rect 33594 46560 33600 46572
rect 33555 46532 33600 46560
rect 33229 46523 33287 46529
rect 33594 46520 33600 46532
rect 33652 46520 33658 46572
rect 34606 46560 34612 46572
rect 34567 46532 34612 46560
rect 34606 46520 34612 46532
rect 34664 46520 34670 46572
rect 35526 46560 35532 46572
rect 35487 46532 35532 46560
rect 35526 46520 35532 46532
rect 35584 46520 35590 46572
rect 36078 46560 36084 46572
rect 36039 46532 36084 46560
rect 36078 46520 36084 46532
rect 36136 46520 36142 46572
rect 37458 46560 37464 46572
rect 37419 46532 37464 46560
rect 37458 46520 37464 46532
rect 37516 46520 37522 46572
rect 37642 46569 37648 46572
rect 37609 46563 37648 46569
rect 37609 46529 37621 46563
rect 37609 46523 37648 46529
rect 37642 46520 37648 46523
rect 37700 46520 37706 46572
rect 37752 46569 37780 46600
rect 40037 46597 40049 46600
rect 40083 46597 40095 46631
rect 40037 46591 40095 46597
rect 40678 46588 40684 46640
rect 40736 46628 40742 46640
rect 41049 46631 41107 46637
rect 41049 46628 41061 46631
rect 40736 46600 41061 46628
rect 40736 46588 40742 46600
rect 41049 46597 41061 46600
rect 41095 46597 41107 46631
rect 41049 46591 41107 46597
rect 37737 46563 37795 46569
rect 37737 46529 37749 46563
rect 37783 46529 37795 46563
rect 37737 46523 37795 46529
rect 33318 46492 33324 46504
rect 33279 46464 33324 46492
rect 33318 46452 33324 46464
rect 33376 46452 33382 46504
rect 33505 46495 33563 46501
rect 33505 46461 33517 46495
rect 33551 46461 33563 46495
rect 33505 46455 33563 46461
rect 32766 46384 32772 46436
rect 32824 46424 32830 46436
rect 33520 46424 33548 46455
rect 33778 46452 33784 46504
rect 33836 46492 33842 46504
rect 35345 46495 35403 46501
rect 35345 46492 35357 46495
rect 33836 46464 35357 46492
rect 33836 46452 33842 46464
rect 35345 46461 35357 46464
rect 35391 46461 35403 46495
rect 35345 46455 35403 46461
rect 35897 46495 35955 46501
rect 35897 46461 35909 46495
rect 35943 46461 35955 46495
rect 37752 46492 37780 46523
rect 37826 46520 37832 46572
rect 37884 46560 37890 46572
rect 38010 46569 38016 46572
rect 37967 46563 38016 46569
rect 37884 46532 37929 46560
rect 37884 46520 37890 46532
rect 37967 46529 37979 46563
rect 38013 46529 38016 46563
rect 37967 46523 38016 46529
rect 38010 46520 38016 46523
rect 38068 46520 38074 46572
rect 38562 46560 38568 46572
rect 38523 46532 38568 46560
rect 38562 46520 38568 46532
rect 38620 46520 38626 46572
rect 38654 46520 38660 46572
rect 38712 46560 38718 46572
rect 38841 46563 38899 46569
rect 38712 46532 38757 46560
rect 38712 46520 38718 46532
rect 38841 46529 38853 46563
rect 38887 46529 38899 46563
rect 38841 46523 38899 46529
rect 38933 46563 38991 46569
rect 38933 46529 38945 46563
rect 38979 46529 38991 46563
rect 38933 46523 38991 46529
rect 38856 46492 38884 46523
rect 37752 46464 38884 46492
rect 38948 46492 38976 46523
rect 39022 46520 39028 46572
rect 39080 46569 39086 46572
rect 39080 46560 39088 46569
rect 39080 46532 39125 46560
rect 39080 46523 39088 46532
rect 39080 46520 39086 46523
rect 39206 46520 39212 46572
rect 39264 46560 39270 46572
rect 39669 46563 39727 46569
rect 39669 46560 39681 46563
rect 39264 46532 39681 46560
rect 39264 46520 39270 46532
rect 39669 46529 39681 46532
rect 39715 46529 39727 46563
rect 39669 46523 39727 46529
rect 39758 46520 39764 46572
rect 39816 46560 39822 46572
rect 39945 46563 40003 46569
rect 39816 46532 39861 46560
rect 39816 46520 39822 46532
rect 39945 46529 39957 46563
rect 39991 46560 40003 46563
rect 40134 46563 40192 46569
rect 39991 46532 40081 46560
rect 39991 46529 40003 46532
rect 39945 46523 40003 46529
rect 39776 46492 39804 46520
rect 38948 46464 39804 46492
rect 35897 46455 35955 46461
rect 35912 46424 35940 46455
rect 38626 46436 38654 46464
rect 36446 46424 36452 46436
rect 32824 46396 36452 46424
rect 32824 46384 32830 46396
rect 36446 46384 36452 46396
rect 36504 46384 36510 46436
rect 37366 46384 37372 46436
rect 37424 46424 37430 46436
rect 37826 46424 37832 46436
rect 37424 46396 37832 46424
rect 37424 46384 37430 46396
rect 37826 46384 37832 46396
rect 37884 46424 37890 46436
rect 38470 46424 38476 46436
rect 37884 46396 38476 46424
rect 37884 46384 37890 46396
rect 38470 46384 38476 46396
rect 38528 46384 38534 46436
rect 38562 46384 38568 46436
rect 38620 46396 38654 46436
rect 40053 46424 40081 46532
rect 40134 46529 40146 46563
rect 40180 46529 40192 46563
rect 40134 46523 40192 46529
rect 40149 46492 40177 46523
rect 40310 46520 40316 46572
rect 40368 46560 40374 46572
rect 41248 46569 41276 46668
rect 41414 46656 41420 46708
rect 41472 46696 41478 46708
rect 43254 46696 43260 46708
rect 41472 46668 41517 46696
rect 43215 46668 43260 46696
rect 41472 46656 41478 46668
rect 43254 46656 43260 46668
rect 43312 46656 43318 46708
rect 44453 46699 44511 46705
rect 43457 46668 44312 46696
rect 42518 46588 42524 46640
rect 42576 46628 42582 46640
rect 42978 46628 42984 46640
rect 42576 46600 42984 46628
rect 42576 46588 42582 46600
rect 42978 46588 42984 46600
rect 43036 46588 43042 46640
rect 40773 46563 40831 46569
rect 40773 46560 40785 46563
rect 40368 46532 40785 46560
rect 40368 46520 40374 46532
rect 40773 46529 40785 46532
rect 40819 46529 40831 46563
rect 40773 46523 40831 46529
rect 40921 46563 40979 46569
rect 40921 46529 40933 46563
rect 40967 46560 40979 46563
rect 41141 46563 41199 46569
rect 40967 46529 41000 46560
rect 40921 46523 41000 46529
rect 41141 46529 41153 46563
rect 41187 46529 41199 46563
rect 41141 46523 41199 46529
rect 41238 46563 41296 46569
rect 41238 46529 41250 46563
rect 41284 46529 41296 46563
rect 41238 46523 41296 46529
rect 40149 46464 40816 46492
rect 40788 46436 40816 46464
rect 40218 46424 40224 46436
rect 40053 46396 40224 46424
rect 38620 46384 38626 46396
rect 40218 46384 40224 46396
rect 40276 46424 40282 46436
rect 40678 46424 40684 46436
rect 40276 46396 40684 46424
rect 40276 46384 40282 46396
rect 40678 46384 40684 46396
rect 40736 46384 40742 46436
rect 40770 46384 40776 46436
rect 40828 46384 40834 46436
rect 40972 46424 41000 46523
rect 41156 46492 41184 46523
rect 42058 46520 42064 46572
rect 42116 46560 42122 46572
rect 42613 46563 42671 46569
rect 42613 46560 42625 46563
rect 42116 46532 42625 46560
rect 42116 46520 42122 46532
rect 42613 46529 42625 46532
rect 42659 46529 42671 46563
rect 42613 46523 42671 46529
rect 42702 46520 42708 46572
rect 42760 46560 42766 46572
rect 42889 46563 42947 46569
rect 42760 46532 42805 46560
rect 42760 46520 42766 46532
rect 42889 46529 42901 46563
rect 42935 46529 42947 46563
rect 43070 46560 43076 46572
rect 43029 46532 43076 46560
rect 42889 46523 42947 46529
rect 41322 46492 41328 46504
rect 41156 46464 41328 46492
rect 41322 46452 41328 46464
rect 41380 46452 41386 46504
rect 42904 46492 42932 46523
rect 43070 46520 43076 46532
rect 43128 46569 43134 46572
rect 43128 46563 43177 46569
rect 43128 46529 43131 46563
rect 43165 46560 43177 46563
rect 43457 46560 43485 46668
rect 43714 46588 43720 46640
rect 43772 46628 43778 46640
rect 44085 46631 44143 46637
rect 44085 46628 44097 46631
rect 43772 46600 44097 46628
rect 43772 46588 43778 46600
rect 44085 46597 44097 46600
rect 44131 46597 44143 46631
rect 44085 46591 44143 46597
rect 44284 46572 44312 46668
rect 44453 46665 44465 46699
rect 44499 46696 44511 46699
rect 45370 46696 45376 46708
rect 44499 46668 45376 46696
rect 44499 46665 44511 46668
rect 44453 46659 44511 46665
rect 45370 46656 45376 46668
rect 45428 46656 45434 46708
rect 46017 46631 46075 46637
rect 46017 46597 46029 46631
rect 46063 46628 46075 46631
rect 46063 46600 48084 46628
rect 46063 46597 46075 46600
rect 46017 46591 46075 46597
rect 43806 46560 43812 46572
rect 43165 46532 43485 46560
rect 43767 46532 43812 46560
rect 43165 46529 43177 46532
rect 43128 46523 43177 46529
rect 43128 46520 43134 46523
rect 43806 46520 43812 46532
rect 43864 46520 43870 46572
rect 43957 46563 44015 46569
rect 43957 46529 43969 46563
rect 44003 46560 44015 46563
rect 44174 46560 44180 46572
rect 44003 46529 44036 46560
rect 44135 46532 44180 46560
rect 43957 46523 44036 46529
rect 43714 46492 43720 46504
rect 42904 46464 43720 46492
rect 43714 46452 43720 46464
rect 43772 46452 43778 46504
rect 41506 46424 41512 46436
rect 40972 46396 41512 46424
rect 41506 46384 41512 46396
rect 41564 46424 41570 46436
rect 41966 46424 41972 46436
rect 41564 46396 41972 46424
rect 41564 46384 41570 46396
rect 41966 46384 41972 46396
rect 42024 46384 42030 46436
rect 44008 46424 44036 46523
rect 44174 46520 44180 46532
rect 44232 46520 44238 46572
rect 44266 46520 44272 46572
rect 44324 46569 44330 46572
rect 44324 46560 44332 46569
rect 45002 46560 45008 46572
rect 44324 46532 44369 46560
rect 44963 46532 45008 46560
rect 44324 46523 44332 46532
rect 44324 46520 44330 46523
rect 45002 46520 45008 46532
rect 45060 46520 45066 46572
rect 45094 46520 45100 46572
rect 45152 46560 45158 46572
rect 45189 46563 45247 46569
rect 45189 46560 45201 46563
rect 45152 46532 45201 46560
rect 45152 46520 45158 46532
rect 45189 46529 45201 46532
rect 45235 46529 45247 46563
rect 47854 46560 47860 46572
rect 47815 46532 47860 46560
rect 45189 46523 45247 46529
rect 47854 46520 47860 46532
rect 47912 46520 47918 46572
rect 48056 46569 48084 46600
rect 48041 46563 48099 46569
rect 48041 46529 48053 46563
rect 48087 46560 48099 46563
rect 48682 46560 48688 46572
rect 48087 46532 48688 46560
rect 48087 46529 48099 46532
rect 48041 46523 48099 46529
rect 48682 46520 48688 46532
rect 48740 46520 48746 46572
rect 48958 46520 48964 46572
rect 49016 46560 49022 46572
rect 49329 46563 49387 46569
rect 49329 46560 49341 46563
rect 49016 46532 49341 46560
rect 49016 46520 49022 46532
rect 49329 46529 49341 46532
rect 49375 46529 49387 46563
rect 49329 46523 49387 46529
rect 48774 46492 48780 46504
rect 48735 46464 48780 46492
rect 48774 46452 48780 46464
rect 48832 46452 48838 46504
rect 49513 46495 49571 46501
rect 49513 46461 49525 46495
rect 49559 46461 49571 46495
rect 49513 46455 49571 46461
rect 44634 46424 44640 46436
rect 44008 46396 44640 46424
rect 31757 46359 31815 46365
rect 31757 46325 31769 46359
rect 31803 46356 31815 46359
rect 31846 46356 31852 46368
rect 31803 46328 31852 46356
rect 31803 46325 31815 46328
rect 31757 46319 31815 46325
rect 31846 46316 31852 46328
rect 31904 46316 31910 46368
rect 32674 46316 32680 46368
rect 32732 46356 32738 46368
rect 33594 46356 33600 46368
rect 32732 46328 33600 46356
rect 32732 46316 32738 46328
rect 33594 46316 33600 46328
rect 33652 46316 33658 46368
rect 38654 46316 38660 46368
rect 38712 46356 38718 46368
rect 41046 46356 41052 46368
rect 38712 46328 41052 46356
rect 38712 46316 38718 46328
rect 41046 46316 41052 46328
rect 41104 46356 41110 46368
rect 41877 46359 41935 46365
rect 41877 46356 41889 46359
rect 41104 46328 41889 46356
rect 41104 46316 41110 46328
rect 41877 46325 41889 46328
rect 41923 46356 41935 46359
rect 44008 46356 44036 46396
rect 44634 46384 44640 46396
rect 44692 46424 44698 46436
rect 48038 46424 48044 46436
rect 44692 46396 48044 46424
rect 44692 46384 44698 46396
rect 48038 46384 48044 46396
rect 48096 46424 48102 46436
rect 49528 46424 49556 46455
rect 48096 46396 49556 46424
rect 48096 46384 48102 46396
rect 41923 46328 44036 46356
rect 41923 46325 41935 46328
rect 41877 46319 41935 46325
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 31754 46112 31760 46164
rect 31812 46152 31818 46164
rect 31812 46124 31857 46152
rect 31812 46112 31818 46124
rect 32490 46112 32496 46164
rect 32548 46152 32554 46164
rect 32953 46155 33011 46161
rect 32953 46152 32965 46155
rect 32548 46124 32965 46152
rect 32548 46112 32554 46124
rect 32953 46121 32965 46124
rect 32999 46121 33011 46155
rect 32953 46115 33011 46121
rect 33689 46155 33747 46161
rect 33689 46121 33701 46155
rect 33735 46152 33747 46155
rect 34606 46152 34612 46164
rect 33735 46124 34612 46152
rect 33735 46121 33747 46124
rect 33689 46115 33747 46121
rect 34606 46112 34612 46124
rect 34664 46112 34670 46164
rect 35526 46112 35532 46164
rect 35584 46152 35590 46164
rect 38286 46152 38292 46164
rect 35584 46124 38292 46152
rect 35584 46112 35590 46124
rect 32582 46044 32588 46096
rect 32640 46084 32646 46096
rect 35342 46084 35348 46096
rect 32640 46056 35348 46084
rect 32640 46044 32646 46056
rect 31021 46019 31079 46025
rect 31021 45985 31033 46019
rect 31067 46016 31079 46019
rect 31067 45988 31616 46016
rect 31067 45985 31079 45988
rect 31021 45979 31079 45985
rect 31478 45948 31484 45960
rect 31439 45920 31484 45948
rect 31478 45908 31484 45920
rect 31536 45908 31542 45960
rect 31588 45957 31616 45988
rect 32674 45976 32680 46028
rect 32732 45976 32738 46028
rect 31573 45951 31631 45957
rect 31573 45917 31585 45951
rect 31619 45948 31631 45951
rect 32122 45948 32128 45960
rect 31619 45920 32128 45948
rect 31619 45917 31631 45920
rect 31573 45911 31631 45917
rect 32122 45908 32128 45920
rect 32180 45908 32186 45960
rect 32306 45948 32312 45960
rect 32267 45920 32312 45948
rect 32306 45908 32312 45920
rect 32364 45908 32370 45960
rect 32457 45951 32515 45957
rect 32457 45917 32469 45951
rect 32503 45948 32515 45951
rect 32692 45948 32720 45976
rect 32784 45957 32812 46056
rect 35342 46044 35348 46056
rect 35400 46044 35406 46096
rect 33318 45976 33324 46028
rect 33376 46016 33382 46028
rect 33376 45988 34192 46016
rect 33376 45976 33382 45988
rect 32503 45920 32720 45948
rect 32774 45951 32832 45957
rect 32503 45917 32515 45920
rect 32457 45911 32515 45917
rect 32774 45917 32786 45951
rect 32820 45917 32832 45951
rect 33410 45948 33416 45960
rect 33371 45920 33416 45948
rect 32774 45911 32832 45917
rect 33410 45908 33416 45920
rect 33468 45908 33474 45960
rect 34164 45957 34192 45988
rect 34238 45976 34244 46028
rect 34296 46016 34302 46028
rect 35544 46016 35572 46112
rect 34296 45988 35572 46016
rect 34296 45976 34302 45988
rect 34149 45951 34207 45957
rect 34149 45917 34161 45951
rect 34195 45948 34207 45951
rect 34790 45948 34796 45960
rect 34195 45920 34796 45948
rect 34195 45917 34207 45920
rect 34149 45911 34207 45917
rect 34790 45908 34796 45920
rect 34848 45908 34854 45960
rect 34882 45908 34888 45960
rect 34940 45948 34946 45960
rect 35253 45951 35311 45957
rect 35253 45948 35265 45951
rect 34940 45920 35265 45948
rect 34940 45908 34946 45920
rect 35253 45917 35265 45920
rect 35299 45917 35311 45951
rect 35253 45911 35311 45917
rect 35805 45951 35863 45957
rect 35805 45917 35817 45951
rect 35851 45948 35863 45951
rect 35894 45948 35900 45960
rect 35851 45920 35900 45948
rect 35851 45917 35863 45920
rect 35805 45911 35863 45917
rect 35894 45908 35900 45920
rect 35952 45908 35958 45960
rect 36096 45957 36124 46124
rect 38286 46112 38292 46124
rect 38344 46112 38350 46164
rect 38470 46112 38476 46164
rect 38528 46152 38534 46164
rect 40494 46152 40500 46164
rect 38528 46124 40500 46152
rect 38528 46112 38534 46124
rect 40494 46112 40500 46124
rect 40552 46152 40558 46164
rect 41049 46155 41107 46161
rect 40552 46124 41000 46152
rect 40552 46112 40558 46124
rect 37642 46044 37648 46096
rect 37700 46084 37706 46096
rect 37700 46056 38608 46084
rect 37700 46044 37706 46056
rect 36173 46019 36231 46025
rect 36173 45985 36185 46019
rect 36219 45985 36231 46019
rect 36446 46016 36452 46028
rect 36407 45988 36452 46016
rect 36173 45979 36231 45985
rect 36081 45951 36139 45957
rect 36081 45917 36093 45951
rect 36127 45917 36139 45951
rect 36188 45948 36216 45979
rect 36446 45976 36452 45988
rect 36504 45976 36510 46028
rect 37734 46016 37740 46028
rect 37695 45988 37740 46016
rect 37734 45976 37740 45988
rect 37792 45976 37798 46028
rect 38580 46025 38608 46056
rect 38746 46044 38752 46096
rect 38804 46084 38810 46096
rect 40972 46084 41000 46124
rect 41049 46121 41061 46155
rect 41095 46152 41107 46155
rect 41230 46152 41236 46164
rect 41095 46124 41236 46152
rect 41095 46121 41107 46124
rect 41049 46115 41107 46121
rect 41230 46112 41236 46124
rect 41288 46112 41294 46164
rect 41966 46152 41972 46164
rect 41879 46124 41972 46152
rect 41966 46112 41972 46124
rect 42024 46152 42030 46164
rect 42702 46152 42708 46164
rect 42024 46124 42708 46152
rect 42024 46112 42030 46124
rect 42702 46112 42708 46124
rect 42760 46112 42766 46164
rect 43162 46112 43168 46164
rect 43220 46152 43226 46164
rect 44174 46152 44180 46164
rect 43220 46124 44180 46152
rect 43220 46112 43226 46124
rect 44174 46112 44180 46124
rect 44232 46112 44238 46164
rect 44269 46155 44327 46161
rect 44269 46121 44281 46155
rect 44315 46152 44327 46155
rect 44450 46152 44456 46164
rect 44315 46124 44456 46152
rect 44315 46121 44327 46124
rect 44269 46115 44327 46121
rect 44450 46112 44456 46124
rect 44508 46112 44514 46164
rect 42518 46084 42524 46096
rect 38804 46056 40908 46084
rect 40972 46056 42524 46084
rect 38804 46044 38810 46056
rect 38565 46019 38623 46025
rect 38565 45985 38577 46019
rect 38611 46016 38623 46019
rect 40880 46016 40908 46056
rect 42518 46044 42524 46056
rect 42576 46044 42582 46096
rect 43990 46084 43996 46096
rect 42904 46056 43996 46084
rect 42904 46025 42932 46056
rect 43990 46044 43996 46056
rect 44048 46044 44054 46096
rect 44192 46084 44220 46112
rect 47026 46084 47032 46096
rect 44192 46056 47032 46084
rect 47026 46044 47032 46056
rect 47084 46044 47090 46096
rect 42889 46019 42947 46025
rect 42889 46016 42901 46019
rect 38611 45988 40816 46016
rect 40880 45988 42901 46016
rect 38611 45985 38623 45988
rect 38565 45979 38623 45985
rect 36354 45948 36360 45960
rect 36188 45920 36360 45948
rect 36081 45911 36139 45917
rect 36354 45908 36360 45920
rect 36412 45908 36418 45960
rect 31757 45883 31815 45889
rect 31757 45849 31769 45883
rect 31803 45880 31815 45883
rect 32140 45880 32168 45908
rect 32585 45883 32643 45889
rect 31803 45852 31892 45880
rect 32140 45852 32444 45880
rect 31803 45849 31815 45852
rect 31757 45843 31815 45849
rect 31864 45824 31892 45852
rect 32416 45824 32444 45852
rect 32585 45849 32597 45883
rect 32631 45849 32643 45883
rect 32585 45843 32643 45849
rect 32677 45883 32735 45889
rect 32677 45849 32689 45883
rect 32723 45880 32735 45883
rect 32950 45880 32956 45892
rect 32723 45852 32956 45880
rect 32723 45849 32735 45852
rect 32677 45843 32735 45849
rect 31846 45772 31852 45824
rect 31904 45772 31910 45824
rect 32398 45772 32404 45824
rect 32456 45772 32462 45824
rect 32600 45812 32628 45843
rect 32950 45840 32956 45852
rect 33008 45840 33014 45892
rect 33686 45880 33692 45892
rect 33599 45852 33692 45880
rect 33686 45840 33692 45852
rect 33744 45880 33750 45892
rect 34330 45880 34336 45892
rect 33744 45852 34336 45880
rect 33744 45840 33750 45852
rect 34330 45840 34336 45852
rect 34388 45840 34394 45892
rect 36464 45880 36492 45976
rect 36722 45948 36728 45960
rect 36683 45920 36728 45948
rect 36722 45908 36728 45920
rect 36780 45908 36786 45960
rect 37550 45948 37556 45960
rect 37511 45920 37556 45948
rect 37550 45908 37556 45920
rect 37608 45908 37614 45960
rect 38286 45908 38292 45960
rect 38344 45948 38350 45960
rect 38381 45951 38439 45957
rect 38381 45948 38393 45951
rect 38344 45920 38393 45948
rect 38344 45908 38350 45920
rect 38381 45917 38393 45920
rect 38427 45917 38439 45951
rect 38838 45948 38844 45960
rect 38799 45920 38844 45948
rect 38381 45911 38439 45917
rect 38838 45908 38844 45920
rect 38896 45908 38902 45960
rect 39209 45951 39267 45957
rect 39209 45917 39221 45951
rect 39255 45917 39267 45951
rect 40402 45948 40408 45960
rect 40363 45920 40408 45948
rect 39209 45911 39267 45917
rect 38654 45880 38660 45892
rect 36464 45852 38660 45880
rect 38654 45840 38660 45852
rect 38712 45880 38718 45892
rect 39224 45880 39252 45911
rect 40402 45908 40408 45920
rect 40460 45908 40466 45960
rect 40494 45908 40500 45960
rect 40552 45948 40558 45960
rect 40552 45920 40597 45948
rect 40552 45908 40558 45920
rect 38712 45852 39252 45880
rect 38712 45840 38718 45852
rect 40218 45840 40224 45892
rect 40276 45880 40282 45892
rect 40788 45889 40816 45988
rect 42889 45985 42901 45988
rect 42935 45985 42947 46019
rect 42889 45979 42947 45985
rect 43070 45976 43076 46028
rect 43128 46016 43134 46028
rect 43128 45988 45324 46016
rect 43128 45976 43134 45988
rect 40862 45908 40868 45960
rect 40920 45957 40926 45960
rect 40920 45948 40928 45957
rect 40920 45920 40965 45948
rect 40920 45911 40928 45920
rect 40920 45908 40926 45911
rect 42518 45908 42524 45960
rect 42576 45948 42582 45960
rect 42613 45951 42671 45957
rect 42613 45948 42625 45951
rect 42576 45920 42625 45948
rect 42576 45908 42582 45920
rect 42613 45917 42625 45920
rect 42659 45917 42671 45951
rect 43622 45948 43628 45960
rect 43583 45920 43628 45948
rect 42613 45911 42671 45917
rect 43622 45908 43628 45920
rect 43680 45908 43686 45960
rect 43773 45951 43831 45957
rect 43773 45917 43785 45951
rect 43819 45948 43831 45951
rect 44008 45948 44036 45988
rect 43819 45920 44036 45948
rect 44131 45951 44189 45957
rect 43819 45917 43831 45920
rect 43773 45911 43831 45917
rect 44131 45917 44143 45951
rect 44177 45948 44189 45951
rect 44266 45948 44272 45960
rect 44177 45920 44272 45948
rect 44177 45917 44189 45920
rect 44131 45911 44189 45917
rect 44266 45908 44272 45920
rect 44324 45908 44330 45960
rect 40681 45883 40739 45889
rect 40681 45880 40693 45883
rect 40276 45852 40693 45880
rect 40276 45840 40282 45852
rect 40681 45849 40693 45852
rect 40727 45849 40739 45883
rect 40681 45843 40739 45849
rect 40773 45883 40831 45889
rect 40773 45849 40785 45883
rect 40819 45849 40831 45883
rect 40773 45843 40831 45849
rect 41693 45883 41751 45889
rect 41693 45849 41705 45883
rect 41739 45880 41751 45883
rect 41782 45880 41788 45892
rect 41739 45852 41788 45880
rect 41739 45849 41751 45852
rect 41693 45843 41751 45849
rect 33042 45812 33048 45824
rect 32600 45784 33048 45812
rect 33042 45772 33048 45784
rect 33100 45772 33106 45824
rect 33505 45815 33563 45821
rect 33505 45781 33517 45815
rect 33551 45812 33563 45815
rect 33778 45812 33784 45824
rect 33551 45784 33784 45812
rect 33551 45781 33563 45784
rect 33505 45775 33563 45781
rect 33778 45772 33784 45784
rect 33836 45772 33842 45824
rect 35342 45772 35348 45824
rect 35400 45812 35406 45824
rect 38010 45812 38016 45824
rect 35400 45784 38016 45812
rect 35400 45772 35406 45784
rect 38010 45772 38016 45784
rect 38068 45812 38074 45824
rect 38746 45812 38752 45824
rect 38068 45784 38752 45812
rect 38068 45772 38074 45784
rect 38746 45772 38752 45784
rect 38804 45812 38810 45824
rect 39022 45812 39028 45824
rect 38804 45784 39028 45812
rect 38804 45772 38810 45784
rect 39022 45772 39028 45784
rect 39080 45772 39086 45824
rect 40788 45812 40816 45843
rect 41782 45840 41788 45852
rect 41840 45840 41846 45892
rect 43901 45883 43959 45889
rect 43901 45880 43913 45883
rect 43732 45852 43913 45880
rect 43732 45824 43760 45852
rect 43901 45849 43913 45852
rect 43947 45849 43959 45883
rect 43901 45843 43959 45849
rect 43993 45883 44051 45889
rect 43993 45849 44005 45883
rect 44039 45880 44051 45883
rect 44634 45880 44640 45892
rect 44039 45852 44640 45880
rect 44039 45849 44051 45852
rect 43993 45843 44051 45849
rect 44634 45840 44640 45852
rect 44692 45840 44698 45892
rect 41966 45812 41972 45824
rect 40788 45784 41972 45812
rect 41966 45772 41972 45784
rect 42024 45772 42030 45824
rect 43714 45772 43720 45824
rect 43772 45772 43778 45824
rect 45296 45821 45324 45988
rect 48498 45948 48504 45960
rect 48459 45920 48504 45948
rect 48498 45908 48504 45920
rect 48556 45908 48562 45960
rect 48682 45948 48688 45960
rect 48643 45920 48688 45948
rect 48682 45908 48688 45920
rect 48740 45908 48746 45960
rect 46198 45880 46204 45892
rect 46159 45852 46204 45880
rect 46198 45840 46204 45852
rect 46256 45880 46262 45892
rect 46845 45883 46903 45889
rect 46845 45880 46857 45883
rect 46256 45852 46857 45880
rect 46256 45840 46262 45852
rect 46845 45849 46857 45852
rect 46891 45880 46903 45883
rect 47118 45880 47124 45892
rect 46891 45852 47124 45880
rect 46891 45849 46903 45852
rect 46845 45843 46903 45849
rect 47118 45840 47124 45852
rect 47176 45840 47182 45892
rect 45281 45815 45339 45821
rect 45281 45781 45293 45815
rect 45327 45812 45339 45815
rect 49326 45812 49332 45824
rect 45327 45784 49332 45812
rect 45327 45781 45339 45784
rect 45281 45775 45339 45781
rect 49326 45772 49332 45784
rect 49384 45772 49390 45824
rect 49510 45812 49516 45824
rect 49471 45784 49516 45812
rect 49510 45772 49516 45784
rect 49568 45772 49574 45824
rect 50433 45815 50491 45821
rect 50433 45781 50445 45815
rect 50479 45812 50491 45815
rect 50798 45812 50804 45824
rect 50479 45784 50804 45812
rect 50479 45781 50491 45784
rect 50433 45775 50491 45781
rect 50798 45772 50804 45784
rect 50856 45772 50862 45824
rect 51629 45815 51687 45821
rect 51629 45781 51641 45815
rect 51675 45812 51687 45815
rect 52086 45812 52092 45824
rect 51675 45784 52092 45812
rect 51675 45781 51687 45784
rect 51629 45775 51687 45781
rect 52086 45772 52092 45784
rect 52144 45772 52150 45824
rect 1104 45722 58880 45744
rect 1104 45670 4874 45722
rect 4926 45670 4938 45722
rect 4990 45670 5002 45722
rect 5054 45670 5066 45722
rect 5118 45670 5130 45722
rect 5182 45670 35594 45722
rect 35646 45670 35658 45722
rect 35710 45670 35722 45722
rect 35774 45670 35786 45722
rect 35838 45670 35850 45722
rect 35902 45670 58880 45722
rect 1104 45648 58880 45670
rect 31846 45608 31852 45620
rect 31128 45580 31852 45608
rect 30561 45475 30619 45481
rect 30561 45441 30573 45475
rect 30607 45472 30619 45475
rect 31021 45475 31079 45481
rect 31021 45472 31033 45475
rect 30607 45444 31033 45472
rect 30607 45441 30619 45444
rect 30561 45435 30619 45441
rect 31021 45441 31033 45444
rect 31067 45472 31079 45475
rect 31128 45472 31156 45580
rect 31846 45568 31852 45580
rect 31904 45608 31910 45620
rect 33686 45608 33692 45620
rect 31904 45580 33692 45608
rect 31904 45568 31910 45580
rect 33686 45568 33692 45580
rect 33744 45568 33750 45620
rect 34241 45611 34299 45617
rect 34241 45577 34253 45611
rect 34287 45608 34299 45611
rect 34514 45608 34520 45620
rect 34287 45580 34520 45608
rect 34287 45577 34299 45580
rect 34241 45571 34299 45577
rect 34514 45568 34520 45580
rect 34572 45608 34578 45620
rect 36354 45608 36360 45620
rect 34572 45580 36360 45608
rect 34572 45568 34578 45580
rect 36354 45568 36360 45580
rect 36412 45568 36418 45620
rect 41877 45611 41935 45617
rect 41877 45577 41889 45611
rect 41923 45608 41935 45611
rect 41966 45608 41972 45620
rect 41923 45580 41972 45608
rect 41923 45577 41935 45580
rect 41877 45571 41935 45577
rect 41966 45568 41972 45580
rect 42024 45568 42030 45620
rect 43441 45611 43499 45617
rect 43441 45577 43453 45611
rect 43487 45608 43499 45611
rect 43622 45608 43628 45620
rect 43487 45580 43628 45608
rect 43487 45577 43499 45580
rect 43441 45571 43499 45577
rect 43622 45568 43628 45580
rect 43680 45568 43686 45620
rect 43990 45568 43996 45620
rect 44048 45608 44054 45620
rect 44085 45611 44143 45617
rect 44085 45608 44097 45611
rect 44048 45580 44097 45608
rect 44048 45568 44054 45580
rect 44085 45577 44097 45580
rect 44131 45577 44143 45611
rect 44085 45571 44143 45577
rect 48317 45611 48375 45617
rect 48317 45577 48329 45611
rect 48363 45608 48375 45611
rect 48498 45608 48504 45620
rect 48363 45580 48504 45608
rect 48363 45577 48375 45580
rect 48317 45571 48375 45577
rect 48498 45568 48504 45580
rect 48556 45568 48562 45620
rect 31570 45500 31576 45552
rect 31628 45540 31634 45552
rect 33410 45540 33416 45552
rect 31628 45512 33416 45540
rect 31628 45500 31634 45512
rect 33410 45500 33416 45512
rect 33468 45540 33474 45552
rect 36725 45543 36783 45549
rect 33468 45512 36676 45540
rect 33468 45500 33474 45512
rect 31067 45444 31156 45472
rect 31205 45475 31263 45481
rect 31067 45441 31079 45444
rect 31021 45435 31079 45441
rect 31205 45441 31217 45475
rect 31251 45441 31263 45475
rect 31205 45435 31263 45441
rect 31297 45475 31355 45481
rect 31297 45441 31309 45475
rect 31343 45472 31355 45475
rect 31588 45472 31616 45500
rect 32398 45472 32404 45484
rect 31343 45444 31616 45472
rect 32359 45444 32404 45472
rect 31343 45441 31355 45444
rect 31297 45435 31355 45441
rect 31220 45404 31248 45435
rect 32398 45432 32404 45444
rect 32456 45432 32462 45484
rect 32769 45475 32827 45481
rect 32769 45441 32781 45475
rect 32815 45472 32827 45475
rect 33318 45472 33324 45484
rect 32815 45444 33324 45472
rect 32815 45441 32827 45444
rect 32769 45435 32827 45441
rect 33318 45432 33324 45444
rect 33376 45432 33382 45484
rect 34164 45481 34192 45512
rect 36648 45484 36676 45512
rect 36725 45509 36737 45543
rect 36771 45540 36783 45543
rect 37642 45540 37648 45552
rect 36771 45512 37648 45540
rect 36771 45509 36783 45512
rect 36725 45503 36783 45509
rect 37642 45500 37648 45512
rect 37700 45500 37706 45552
rect 39853 45543 39911 45549
rect 39853 45509 39865 45543
rect 39899 45509 39911 45543
rect 39853 45503 39911 45509
rect 34149 45475 34207 45481
rect 34149 45441 34161 45475
rect 34195 45441 34207 45475
rect 34149 45435 34207 45441
rect 34330 45432 34336 45484
rect 34388 45472 34394 45484
rect 34425 45475 34483 45481
rect 34425 45472 34437 45475
rect 34388 45444 34437 45472
rect 34388 45432 34394 45444
rect 34425 45441 34437 45444
rect 34471 45441 34483 45475
rect 34425 45435 34483 45441
rect 35069 45475 35127 45481
rect 35069 45441 35081 45475
rect 35115 45472 35127 45475
rect 35434 45472 35440 45484
rect 35115 45444 35440 45472
rect 35115 45441 35127 45444
rect 35069 45435 35127 45441
rect 35434 45432 35440 45444
rect 35492 45432 35498 45484
rect 36630 45472 36636 45484
rect 36591 45444 36636 45472
rect 36630 45432 36636 45444
rect 36688 45432 36694 45484
rect 36909 45475 36967 45481
rect 36909 45441 36921 45475
rect 36955 45472 36967 45475
rect 37458 45472 37464 45484
rect 36955 45444 37464 45472
rect 36955 45441 36967 45444
rect 36909 45435 36967 45441
rect 31846 45404 31852 45416
rect 31220 45376 31852 45404
rect 31846 45364 31852 45376
rect 31904 45364 31910 45416
rect 34514 45364 34520 45416
rect 34572 45404 34578 45416
rect 34977 45407 35035 45413
rect 34977 45404 34989 45407
rect 34572 45376 34989 45404
rect 34572 45364 34578 45376
rect 34977 45373 34989 45376
rect 35023 45373 35035 45407
rect 36924 45404 36952 45435
rect 37458 45432 37464 45444
rect 37516 45432 37522 45484
rect 37734 45432 37740 45484
rect 37792 45472 37798 45484
rect 38197 45475 38255 45481
rect 38197 45472 38209 45475
rect 37792 45444 38209 45472
rect 37792 45432 37798 45444
rect 38197 45441 38209 45444
rect 38243 45441 38255 45475
rect 38197 45435 38255 45441
rect 39206 45432 39212 45484
rect 39264 45472 39270 45484
rect 39577 45475 39635 45481
rect 39577 45472 39589 45475
rect 39264 45444 39589 45472
rect 39264 45432 39270 45444
rect 39577 45441 39589 45444
rect 39623 45441 39635 45475
rect 39868 45472 39896 45503
rect 40218 45500 40224 45552
rect 40276 45540 40282 45552
rect 40589 45543 40647 45549
rect 40589 45540 40601 45543
rect 40276 45512 40601 45540
rect 40276 45500 40282 45512
rect 40589 45509 40601 45512
rect 40635 45509 40647 45543
rect 41414 45540 41420 45552
rect 40589 45503 40647 45509
rect 40696 45512 41420 45540
rect 40494 45481 40500 45484
rect 40313 45475 40371 45481
rect 40313 45472 40325 45475
rect 39868 45444 40325 45472
rect 39577 45435 39635 45441
rect 40313 45441 40325 45444
rect 40359 45441 40371 45475
rect 40313 45435 40371 45441
rect 40461 45475 40500 45481
rect 40461 45441 40473 45475
rect 40461 45435 40500 45441
rect 40494 45432 40500 45435
rect 40552 45432 40558 45484
rect 40696 45481 40724 45512
rect 41414 45500 41420 45512
rect 41472 45500 41478 45552
rect 43456 45512 44220 45540
rect 40681 45475 40739 45481
rect 40681 45441 40693 45475
rect 40727 45441 40739 45475
rect 40681 45435 40739 45441
rect 34977 45367 35035 45373
rect 36372 45376 36952 45404
rect 34425 45339 34483 45345
rect 34425 45305 34437 45339
rect 34471 45336 34483 45339
rect 34882 45336 34888 45348
rect 34471 45308 34888 45336
rect 34471 45305 34483 45308
rect 34425 45299 34483 45305
rect 34882 45296 34888 45308
rect 34940 45296 34946 45348
rect 35989 45339 36047 45345
rect 35989 45305 36001 45339
rect 36035 45336 36047 45339
rect 36170 45336 36176 45348
rect 36035 45308 36176 45336
rect 36035 45305 36047 45308
rect 35989 45299 36047 45305
rect 36170 45296 36176 45308
rect 36228 45336 36234 45348
rect 36372 45336 36400 45376
rect 37826 45364 37832 45416
rect 37884 45404 37890 45416
rect 38105 45407 38163 45413
rect 38105 45404 38117 45407
rect 37884 45376 38117 45404
rect 37884 45364 37890 45376
rect 38105 45373 38117 45376
rect 38151 45373 38163 45407
rect 38105 45367 38163 45373
rect 39758 45364 39764 45416
rect 39816 45404 39822 45416
rect 39853 45407 39911 45413
rect 39853 45404 39865 45407
rect 39816 45376 39865 45404
rect 39816 45364 39822 45376
rect 39853 45373 39865 45376
rect 39899 45373 39911 45407
rect 39853 45367 39911 45373
rect 36228 45308 36400 45336
rect 36909 45339 36967 45345
rect 36228 45296 36234 45308
rect 36909 45305 36921 45339
rect 36955 45336 36967 45339
rect 37550 45336 37556 45348
rect 36955 45308 37556 45336
rect 36955 45305 36967 45308
rect 36909 45299 36967 45305
rect 37550 45296 37556 45308
rect 37608 45296 37614 45348
rect 39025 45339 39083 45345
rect 39025 45336 39037 45339
rect 37660 45308 39037 45336
rect 31021 45271 31079 45277
rect 31021 45237 31033 45271
rect 31067 45268 31079 45271
rect 31110 45268 31116 45280
rect 31067 45240 31116 45268
rect 31067 45237 31079 45240
rect 31021 45231 31079 45237
rect 31110 45228 31116 45240
rect 31168 45228 31174 45280
rect 35342 45268 35348 45280
rect 35303 45240 35348 45268
rect 35342 45228 35348 45240
rect 35400 45228 35406 45280
rect 37458 45268 37464 45280
rect 37419 45240 37464 45268
rect 37458 45228 37464 45240
rect 37516 45268 37522 45280
rect 37660 45268 37688 45308
rect 39025 45305 39037 45308
rect 39071 45305 39083 45339
rect 39025 45299 39083 45305
rect 39206 45296 39212 45348
rect 39264 45336 39270 45348
rect 40696 45336 40724 45435
rect 40770 45432 40776 45484
rect 40828 45481 40834 45484
rect 40828 45472 40836 45481
rect 41785 45475 41843 45481
rect 40828 45444 40873 45472
rect 40828 45435 40836 45444
rect 41785 45441 41797 45475
rect 41831 45441 41843 45475
rect 41785 45435 41843 45441
rect 42061 45475 42119 45481
rect 42061 45441 42073 45475
rect 42107 45472 42119 45475
rect 42794 45472 42800 45484
rect 42107 45444 42800 45472
rect 42107 45441 42119 45444
rect 42061 45435 42119 45441
rect 40828 45432 40834 45435
rect 41800 45404 41828 45435
rect 42794 45432 42800 45444
rect 42852 45432 42858 45484
rect 43162 45472 43168 45484
rect 43123 45444 43168 45472
rect 43162 45432 43168 45444
rect 43220 45432 43226 45484
rect 42886 45404 42892 45416
rect 41800 45376 42892 45404
rect 42886 45364 42892 45376
rect 42944 45404 42950 45416
rect 43456 45413 43484 45512
rect 44192 45481 44220 45512
rect 47026 45500 47032 45552
rect 47084 45540 47090 45552
rect 47084 45512 49372 45540
rect 47084 45500 47090 45512
rect 43901 45475 43959 45481
rect 43901 45472 43913 45475
rect 43732 45444 43913 45472
rect 43441 45407 43499 45413
rect 43441 45404 43453 45407
rect 42944 45376 43453 45404
rect 42944 45364 42950 45376
rect 43441 45373 43453 45376
rect 43487 45373 43499 45407
rect 43441 45367 43499 45373
rect 40954 45336 40960 45348
rect 39264 45308 40724 45336
rect 40915 45308 40960 45336
rect 39264 45296 39270 45308
rect 40954 45296 40960 45308
rect 41012 45296 41018 45348
rect 42058 45336 42064 45348
rect 42019 45308 42064 45336
rect 42058 45296 42064 45308
rect 42116 45296 42122 45348
rect 42705 45339 42763 45345
rect 42705 45305 42717 45339
rect 42751 45336 42763 45339
rect 43070 45336 43076 45348
rect 42751 45308 43076 45336
rect 42751 45305 42763 45308
rect 42705 45299 42763 45305
rect 37516 45240 37688 45268
rect 38473 45271 38531 45277
rect 37516 45228 37522 45240
rect 38473 45237 38485 45271
rect 38519 45268 38531 45271
rect 38930 45268 38936 45280
rect 38519 45240 38936 45268
rect 38519 45237 38531 45240
rect 38473 45231 38531 45237
rect 38930 45228 38936 45240
rect 38988 45228 38994 45280
rect 39298 45228 39304 45280
rect 39356 45268 39362 45280
rect 39669 45271 39727 45277
rect 39669 45268 39681 45271
rect 39356 45240 39681 45268
rect 39356 45228 39362 45240
rect 39669 45237 39681 45240
rect 39715 45237 39727 45271
rect 39669 45231 39727 45237
rect 41414 45228 41420 45280
rect 41472 45268 41478 45280
rect 42720 45268 42748 45299
rect 43070 45296 43076 45308
rect 43128 45296 43134 45348
rect 43732 45336 43760 45444
rect 43901 45441 43913 45444
rect 43947 45441 43959 45475
rect 43901 45435 43959 45441
rect 44177 45475 44235 45481
rect 44177 45441 44189 45475
rect 44223 45441 44235 45475
rect 45002 45472 45008 45484
rect 44963 45444 45008 45472
rect 44177 45435 44235 45441
rect 45002 45432 45008 45444
rect 45060 45432 45066 45484
rect 45094 45432 45100 45484
rect 45152 45472 45158 45484
rect 49344 45481 49372 45512
rect 46293 45475 46351 45481
rect 46293 45472 46305 45475
rect 45152 45444 46305 45472
rect 45152 45432 45158 45444
rect 46293 45441 46305 45444
rect 46339 45441 46351 45475
rect 46293 45435 46351 45441
rect 47949 45475 48007 45481
rect 47949 45441 47961 45475
rect 47995 45441 48007 45475
rect 47949 45435 48007 45441
rect 49329 45475 49387 45481
rect 49329 45441 49341 45475
rect 49375 45441 49387 45475
rect 49329 45435 49387 45441
rect 43806 45364 43812 45416
rect 43864 45404 43870 45416
rect 44913 45407 44971 45413
rect 44913 45404 44925 45407
rect 43864 45376 44925 45404
rect 43864 45364 43870 45376
rect 44913 45373 44925 45376
rect 44959 45373 44971 45407
rect 44913 45367 44971 45373
rect 45738 45364 45744 45416
rect 45796 45404 45802 45416
rect 46201 45407 46259 45413
rect 46201 45404 46213 45407
rect 45796 45376 46213 45404
rect 45796 45364 45802 45376
rect 46201 45373 46213 45376
rect 46247 45373 46259 45407
rect 46201 45367 46259 45373
rect 47964 45348 47992 45435
rect 49418 45432 49424 45484
rect 49476 45472 49482 45484
rect 50709 45475 50767 45481
rect 50709 45472 50721 45475
rect 49476 45444 50721 45472
rect 49476 45432 49482 45444
rect 50709 45441 50721 45444
rect 50755 45441 50767 45475
rect 50709 45435 50767 45441
rect 48041 45407 48099 45413
rect 48041 45373 48053 45407
rect 48087 45404 48099 45407
rect 48406 45404 48412 45416
rect 48087 45376 48412 45404
rect 48087 45373 48099 45376
rect 48041 45367 48099 45373
rect 48406 45364 48412 45376
rect 48464 45364 48470 45416
rect 49513 45407 49571 45413
rect 49513 45373 49525 45407
rect 49559 45373 49571 45407
rect 50890 45404 50896 45416
rect 50851 45376 50896 45404
rect 49513 45367 49571 45373
rect 43898 45336 43904 45348
rect 43272 45308 43760 45336
rect 43859 45308 43904 45336
rect 41472 45240 42748 45268
rect 41472 45228 41478 45240
rect 42794 45228 42800 45280
rect 42852 45268 42858 45280
rect 43272 45277 43300 45308
rect 43898 45296 43904 45308
rect 43956 45296 43962 45348
rect 45373 45339 45431 45345
rect 45373 45305 45385 45339
rect 45419 45336 45431 45339
rect 47946 45336 47952 45348
rect 45419 45308 47952 45336
rect 45419 45305 45431 45308
rect 45373 45299 45431 45305
rect 47946 45296 47952 45308
rect 48004 45296 48010 45348
rect 49326 45296 49332 45348
rect 49384 45336 49390 45348
rect 49528 45336 49556 45367
rect 50890 45364 50896 45376
rect 50948 45364 50954 45416
rect 51534 45404 51540 45416
rect 51495 45376 51540 45404
rect 51534 45364 51540 45376
rect 51592 45364 51598 45416
rect 49384 45308 49556 45336
rect 49384 45296 49390 45308
rect 50798 45296 50804 45348
rect 50856 45336 50862 45348
rect 51997 45339 52055 45345
rect 51997 45336 52009 45339
rect 50856 45308 52009 45336
rect 50856 45296 50862 45308
rect 51997 45305 52009 45308
rect 52043 45305 52055 45339
rect 51997 45299 52055 45305
rect 43257 45271 43315 45277
rect 43257 45268 43269 45271
rect 42852 45240 43269 45268
rect 42852 45228 42858 45240
rect 43257 45237 43269 45240
rect 43303 45237 43315 45271
rect 43257 45231 43315 45237
rect 46569 45271 46627 45277
rect 46569 45237 46581 45271
rect 46615 45268 46627 45271
rect 50522 45268 50528 45280
rect 46615 45240 50528 45268
rect 46615 45237 46627 45240
rect 46569 45231 46627 45237
rect 50522 45228 50528 45240
rect 50580 45228 50586 45280
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 34054 45064 34060 45076
rect 34015 45036 34060 45064
rect 34054 45024 34060 45036
rect 34112 45024 34118 45076
rect 38286 45024 38292 45076
rect 38344 45064 38350 45076
rect 40037 45067 40095 45073
rect 40037 45064 40049 45067
rect 38344 45036 40049 45064
rect 38344 45024 38350 45036
rect 40037 45033 40049 45036
rect 40083 45033 40095 45067
rect 40037 45027 40095 45033
rect 40681 45067 40739 45073
rect 40681 45033 40693 45067
rect 40727 45064 40739 45067
rect 41046 45064 41052 45076
rect 40727 45036 41052 45064
rect 40727 45033 40739 45036
rect 40681 45027 40739 45033
rect 34238 44996 34244 45008
rect 32140 44968 34244 44996
rect 31846 44928 31852 44940
rect 31807 44900 31852 44928
rect 31846 44888 31852 44900
rect 31904 44888 31910 44940
rect 31110 44860 31116 44872
rect 31071 44832 31116 44860
rect 31110 44820 31116 44832
rect 31168 44820 31174 44872
rect 31662 44860 31668 44872
rect 31623 44832 31668 44860
rect 31662 44820 31668 44832
rect 31720 44820 31726 44872
rect 32033 44863 32091 44869
rect 32033 44829 32045 44863
rect 32079 44860 32091 44863
rect 32140 44860 32168 44968
rect 34238 44956 34244 44968
rect 34296 44956 34302 45008
rect 34330 44956 34336 45008
rect 34388 44996 34394 45008
rect 36078 44996 36084 45008
rect 34388 44968 36084 44996
rect 34388 44956 34394 44968
rect 36078 44956 36084 44968
rect 36136 44956 36142 45008
rect 40696 44996 40724 45027
rect 41046 45024 41052 45036
rect 41104 45024 41110 45076
rect 43162 45064 43168 45076
rect 41253 45036 43168 45064
rect 38028 44968 40724 44996
rect 38028 44940 38056 44968
rect 32398 44888 32404 44940
rect 32456 44928 32462 44940
rect 34606 44928 34612 44940
rect 32456 44900 34612 44928
rect 32456 44888 32462 44900
rect 32600 44869 32628 44900
rect 34606 44888 34612 44900
rect 34664 44888 34670 44940
rect 35342 44888 35348 44940
rect 35400 44928 35406 44940
rect 35713 44931 35771 44937
rect 35713 44928 35725 44931
rect 35400 44900 35725 44928
rect 35400 44888 35406 44900
rect 35713 44897 35725 44900
rect 35759 44897 35771 44931
rect 38010 44928 38016 44940
rect 37971 44900 38016 44928
rect 35713 44891 35771 44897
rect 38010 44888 38016 44900
rect 38068 44888 38074 44940
rect 38286 44928 38292 44940
rect 38120 44900 38292 44928
rect 32079 44832 32168 44860
rect 32585 44863 32643 44869
rect 32079 44829 32091 44832
rect 32033 44823 32091 44829
rect 32585 44829 32597 44863
rect 32631 44829 32643 44863
rect 32766 44860 32772 44872
rect 32727 44832 32772 44860
rect 32585 44823 32643 44829
rect 32766 44820 32772 44832
rect 32824 44820 32830 44872
rect 32858 44820 32864 44872
rect 32916 44860 32922 44872
rect 33413 44863 33471 44869
rect 33413 44860 33425 44863
rect 32916 44832 33425 44860
rect 32916 44820 32922 44832
rect 33413 44829 33425 44832
rect 33459 44829 33471 44863
rect 33413 44823 33471 44829
rect 33502 44820 33508 44872
rect 33560 44860 33566 44872
rect 33878 44863 33936 44869
rect 33560 44832 33605 44860
rect 33560 44820 33566 44832
rect 33878 44829 33890 44863
rect 33924 44860 33936 44863
rect 33924 44832 34008 44860
rect 33924 44829 33936 44832
rect 33878 44823 33936 44829
rect 33042 44752 33048 44804
rect 33100 44792 33106 44804
rect 33689 44795 33747 44801
rect 33689 44792 33701 44795
rect 33100 44764 33701 44792
rect 33100 44752 33106 44764
rect 33689 44761 33701 44764
rect 33735 44761 33747 44795
rect 33689 44755 33747 44761
rect 33778 44752 33784 44804
rect 33836 44792 33842 44804
rect 33836 44764 33881 44792
rect 33836 44752 33842 44764
rect 32490 44684 32496 44736
rect 32548 44724 32554 44736
rect 33980 44724 34008 44832
rect 34514 44820 34520 44872
rect 34572 44860 34578 44872
rect 35526 44860 35532 44872
rect 34572 44832 35532 44860
rect 34572 44820 34578 44832
rect 35526 44820 35532 44832
rect 35584 44860 35590 44872
rect 35897 44863 35955 44869
rect 35897 44860 35909 44863
rect 35584 44832 35909 44860
rect 35584 44820 35590 44832
rect 35897 44829 35909 44832
rect 35943 44829 35955 44863
rect 35897 44823 35955 44829
rect 36906 44820 36912 44872
rect 36964 44860 36970 44872
rect 37277 44863 37335 44869
rect 37277 44860 37289 44863
rect 36964 44832 37289 44860
rect 36964 44820 36970 44832
rect 37277 44829 37289 44832
rect 37323 44829 37335 44863
rect 37826 44860 37832 44872
rect 37787 44832 37832 44860
rect 37277 44823 37335 44829
rect 37826 44820 37832 44832
rect 37884 44820 37890 44872
rect 38120 44869 38148 44900
rect 38286 44888 38292 44900
rect 38344 44888 38350 44940
rect 38654 44928 38660 44940
rect 38615 44900 38660 44928
rect 38654 44888 38660 44900
rect 38712 44888 38718 44940
rect 41253 44928 41281 45036
rect 43162 45024 43168 45036
rect 43220 45024 43226 45076
rect 43806 45064 43812 45076
rect 43767 45036 43812 45064
rect 43806 45024 43812 45036
rect 43864 45024 43870 45076
rect 47118 45064 47124 45076
rect 47079 45036 47124 45064
rect 47118 45024 47124 45036
rect 47176 45024 47182 45076
rect 50890 45064 50896 45076
rect 50851 45036 50896 45064
rect 50890 45024 50896 45036
rect 50948 45024 50954 45076
rect 42797 44999 42855 45005
rect 42797 44965 42809 44999
rect 42843 44996 42855 44999
rect 45094 44996 45100 45008
rect 42843 44968 45100 44996
rect 42843 44965 42855 44968
rect 42797 44959 42855 44965
rect 45094 44956 45100 44968
rect 45152 44956 45158 45008
rect 43346 44928 43352 44940
rect 38764 44900 41281 44928
rect 41524 44900 43208 44928
rect 43307 44900 43352 44928
rect 38105 44863 38163 44869
rect 38105 44829 38117 44863
rect 38151 44829 38163 44863
rect 38105 44823 38163 44829
rect 38194 44820 38200 44872
rect 38252 44860 38258 44872
rect 38764 44869 38792 44900
rect 38749 44863 38807 44869
rect 38749 44860 38761 44863
rect 38252 44832 38761 44860
rect 38252 44820 38258 44832
rect 38749 44829 38761 44832
rect 38795 44829 38807 44863
rect 38749 44823 38807 44829
rect 36633 44795 36691 44801
rect 36633 44761 36645 44795
rect 36679 44792 36691 44795
rect 41524 44792 41552 44900
rect 41601 44863 41659 44869
rect 41601 44829 41613 44863
rect 41647 44860 41659 44863
rect 41966 44860 41972 44872
rect 41647 44832 41972 44860
rect 41647 44829 41659 44832
rect 41601 44823 41659 44829
rect 41966 44820 41972 44832
rect 42024 44820 42030 44872
rect 42150 44860 42156 44872
rect 42111 44832 42156 44860
rect 42150 44820 42156 44832
rect 42208 44820 42214 44872
rect 42242 44820 42248 44872
rect 42300 44860 42306 44872
rect 42300 44832 42345 44860
rect 42300 44820 42306 44832
rect 42426 44820 42432 44872
rect 42484 44860 42490 44872
rect 42659 44863 42717 44869
rect 42484 44832 42529 44860
rect 42484 44820 42490 44832
rect 42659 44829 42671 44863
rect 42705 44860 42717 44863
rect 42978 44860 42984 44872
rect 42705 44832 42984 44860
rect 42705 44829 42717 44832
rect 42659 44823 42717 44829
rect 42978 44820 42984 44832
rect 43036 44820 43042 44872
rect 36679 44764 41552 44792
rect 36679 44761 36691 44764
rect 36633 44755 36691 44761
rect 42334 44752 42340 44804
rect 42392 44792 42398 44804
rect 42521 44795 42579 44801
rect 42521 44792 42533 44795
rect 42392 44764 42533 44792
rect 42392 44752 42398 44764
rect 42521 44761 42533 44764
rect 42567 44761 42579 44795
rect 43180 44792 43208 44900
rect 43346 44888 43352 44900
rect 43404 44888 43410 44940
rect 46293 44931 46351 44937
rect 46293 44897 46305 44931
rect 46339 44928 46351 44931
rect 48501 44931 48559 44937
rect 48501 44928 48513 44931
rect 46339 44900 48513 44928
rect 46339 44897 46351 44900
rect 46293 44891 46351 44897
rect 48501 44897 48513 44900
rect 48547 44928 48559 44931
rect 49418 44928 49424 44940
rect 48547 44900 49424 44928
rect 48547 44897 48559 44900
rect 48501 44891 48559 44897
rect 49418 44888 49424 44900
rect 49476 44888 49482 44940
rect 50614 44928 50620 44940
rect 50575 44900 50620 44928
rect 50614 44888 50620 44900
rect 50672 44888 50678 44940
rect 51994 44928 52000 44940
rect 51955 44900 52000 44928
rect 51994 44888 52000 44900
rect 52052 44888 52058 44940
rect 52273 44931 52331 44937
rect 52273 44897 52285 44931
rect 52319 44928 52331 44931
rect 53006 44928 53012 44940
rect 52319 44900 53012 44928
rect 52319 44897 52331 44900
rect 52273 44891 52331 44897
rect 53006 44888 53012 44900
rect 53064 44888 53070 44940
rect 43438 44860 43444 44872
rect 43399 44832 43444 44860
rect 43438 44820 43444 44832
rect 43496 44820 43502 44872
rect 43990 44820 43996 44872
rect 44048 44860 44054 44872
rect 45281 44863 45339 44869
rect 45281 44860 45293 44863
rect 44048 44832 45293 44860
rect 44048 44820 44054 44832
rect 45281 44829 45293 44832
rect 45327 44829 45339 44863
rect 45281 44823 45339 44829
rect 45370 44820 45376 44872
rect 45428 44860 45434 44872
rect 45465 44863 45523 44869
rect 45465 44860 45477 44863
rect 45428 44832 45477 44860
rect 45428 44820 45434 44832
rect 45465 44829 45477 44832
rect 45511 44829 45523 44863
rect 45465 44823 45523 44829
rect 47946 44820 47952 44872
rect 48004 44860 48010 44872
rect 48409 44863 48467 44869
rect 48409 44860 48421 44863
rect 48004 44832 48421 44860
rect 48004 44820 48010 44832
rect 48409 44829 48421 44832
rect 48455 44829 48467 44863
rect 50522 44860 50528 44872
rect 50483 44832 50528 44860
rect 48409 44823 48467 44829
rect 50522 44820 50528 44832
rect 50580 44860 50586 44872
rect 51905 44863 51963 44869
rect 51905 44860 51917 44863
rect 50580 44832 51917 44860
rect 50580 44820 50586 44832
rect 51905 44829 51917 44832
rect 51951 44829 51963 44863
rect 51905 44823 51963 44829
rect 45002 44792 45008 44804
rect 43180 44764 45008 44792
rect 42521 44755 42579 44761
rect 45002 44752 45008 44764
rect 45060 44752 45066 44804
rect 32548 44696 34008 44724
rect 32548 44684 32554 44696
rect 34606 44684 34612 44736
rect 34664 44724 34670 44736
rect 34885 44727 34943 44733
rect 34885 44724 34897 44727
rect 34664 44696 34897 44724
rect 34664 44684 34670 44696
rect 34885 44693 34897 44696
rect 34931 44693 34943 44727
rect 34885 44687 34943 44693
rect 41230 44684 41236 44736
rect 41288 44724 41294 44736
rect 41325 44727 41383 44733
rect 41325 44724 41337 44727
rect 41288 44696 41337 44724
rect 41288 44684 41294 44696
rect 41325 44693 41337 44696
rect 41371 44693 41383 44727
rect 41325 44687 41383 44693
rect 42426 44684 42432 44736
rect 42484 44724 42490 44736
rect 43622 44724 43628 44736
rect 42484 44696 43628 44724
rect 42484 44684 42490 44696
rect 43622 44684 43628 44696
rect 43680 44684 43686 44736
rect 44361 44727 44419 44733
rect 44361 44693 44373 44727
rect 44407 44724 44419 44727
rect 44450 44724 44456 44736
rect 44407 44696 44456 44724
rect 44407 44693 44419 44696
rect 44361 44687 44419 44693
rect 44450 44684 44456 44696
rect 44508 44684 44514 44736
rect 47670 44724 47676 44736
rect 47631 44696 47676 44724
rect 47670 44684 47676 44696
rect 47728 44684 47734 44736
rect 48777 44727 48835 44733
rect 48777 44693 48789 44727
rect 48823 44724 48835 44727
rect 49142 44724 49148 44736
rect 48823 44696 49148 44724
rect 48823 44693 48835 44696
rect 48777 44687 48835 44693
rect 49142 44684 49148 44696
rect 49200 44684 49206 44736
rect 49234 44684 49240 44736
rect 49292 44724 49298 44736
rect 49329 44727 49387 44733
rect 49329 44724 49341 44727
rect 49292 44696 49341 44724
rect 49292 44684 49298 44696
rect 49329 44693 49341 44696
rect 49375 44724 49387 44727
rect 50522 44724 50528 44736
rect 49375 44696 50528 44724
rect 49375 44693 49387 44696
rect 49329 44687 49387 44693
rect 50522 44684 50528 44696
rect 50580 44684 50586 44736
rect 52638 44684 52644 44736
rect 52696 44724 52702 44736
rect 52917 44727 52975 44733
rect 52917 44724 52929 44727
rect 52696 44696 52929 44724
rect 52696 44684 52702 44696
rect 52917 44693 52929 44696
rect 52963 44693 52975 44727
rect 52917 44687 52975 44693
rect 1104 44634 58880 44656
rect 1104 44582 4874 44634
rect 4926 44582 4938 44634
rect 4990 44582 5002 44634
rect 5054 44582 5066 44634
rect 5118 44582 5130 44634
rect 5182 44582 35594 44634
rect 35646 44582 35658 44634
rect 35710 44582 35722 44634
rect 35774 44582 35786 44634
rect 35838 44582 35850 44634
rect 35902 44582 58880 44634
rect 1104 44560 58880 44582
rect 32858 44520 32864 44532
rect 32819 44492 32864 44520
rect 32858 44480 32864 44492
rect 32916 44480 32922 44532
rect 34425 44523 34483 44529
rect 34425 44489 34437 44523
rect 34471 44520 34483 44523
rect 34514 44520 34520 44532
rect 34471 44492 34520 44520
rect 34471 44489 34483 44492
rect 34425 44483 34483 44489
rect 34514 44480 34520 44492
rect 34572 44480 34578 44532
rect 36725 44523 36783 44529
rect 36725 44489 36737 44523
rect 36771 44520 36783 44523
rect 38838 44520 38844 44532
rect 36771 44492 38844 44520
rect 36771 44489 36783 44492
rect 36725 44483 36783 44489
rect 38838 44480 38844 44492
rect 38896 44480 38902 44532
rect 41414 44480 41420 44532
rect 41472 44520 41478 44532
rect 42061 44523 42119 44529
rect 41472 44492 41517 44520
rect 41472 44480 41478 44492
rect 42061 44489 42073 44523
rect 42107 44520 42119 44523
rect 42242 44520 42248 44532
rect 42107 44492 42248 44520
rect 42107 44489 42119 44492
rect 42061 44483 42119 44489
rect 42242 44480 42248 44492
rect 42300 44520 42306 44532
rect 42797 44523 42855 44529
rect 42797 44520 42809 44523
rect 42300 44492 42809 44520
rect 42300 44480 42306 44492
rect 42797 44489 42809 44492
rect 42843 44520 42855 44523
rect 42843 44492 43760 44520
rect 42843 44489 42855 44492
rect 42797 44483 42855 44489
rect 35989 44455 36047 44461
rect 35989 44421 36001 44455
rect 36035 44452 36047 44455
rect 43346 44452 43352 44464
rect 36035 44424 43352 44452
rect 36035 44421 36047 44424
rect 35989 44415 36047 44421
rect 43346 44412 43352 44424
rect 43404 44452 43410 44464
rect 43732 44452 43760 44492
rect 43898 44480 43904 44532
rect 43956 44520 43962 44532
rect 47029 44523 47087 44529
rect 47029 44520 47041 44523
rect 43956 44492 47041 44520
rect 43956 44480 43962 44492
rect 47029 44489 47041 44492
rect 47075 44520 47087 44523
rect 48406 44520 48412 44532
rect 47075 44492 48176 44520
rect 48367 44492 48412 44520
rect 47075 44489 47087 44492
rect 47029 44483 47087 44489
rect 44450 44452 44456 44464
rect 43404 44424 43668 44452
rect 43732 44424 44456 44452
rect 43404 44412 43410 44424
rect 31205 44387 31263 44393
rect 31205 44353 31217 44387
rect 31251 44384 31263 44387
rect 31662 44384 31668 44396
rect 31251 44356 31668 44384
rect 31251 44353 31263 44356
rect 31205 44347 31263 44353
rect 31662 44344 31668 44356
rect 31720 44344 31726 44396
rect 32585 44387 32643 44393
rect 32585 44353 32597 44387
rect 32631 44384 32643 44387
rect 33318 44384 33324 44396
rect 32631 44356 33324 44384
rect 32631 44353 32643 44356
rect 32585 44347 32643 44353
rect 33318 44344 33324 44356
rect 33376 44344 33382 44396
rect 33781 44387 33839 44393
rect 33781 44353 33793 44387
rect 33827 44384 33839 44387
rect 34054 44384 34060 44396
rect 33827 44356 34060 44384
rect 33827 44353 33839 44356
rect 33781 44347 33839 44353
rect 34054 44344 34060 44356
rect 34112 44344 34118 44396
rect 34514 44344 34520 44396
rect 34572 44384 34578 44396
rect 34977 44387 35035 44393
rect 34977 44384 34989 44387
rect 34572 44356 34989 44384
rect 34572 44344 34578 44356
rect 34977 44353 34989 44356
rect 35023 44353 35035 44387
rect 34977 44347 35035 44353
rect 35161 44387 35219 44393
rect 35161 44353 35173 44387
rect 35207 44353 35219 44387
rect 36630 44384 36636 44396
rect 36543 44356 36636 44384
rect 35161 44347 35219 44353
rect 31018 44276 31024 44328
rect 31076 44316 31082 44328
rect 31113 44319 31171 44325
rect 31113 44316 31125 44319
rect 31076 44288 31125 44316
rect 31076 44276 31082 44288
rect 31113 44285 31125 44288
rect 31159 44285 31171 44319
rect 31113 44279 31171 44285
rect 32398 44276 32404 44328
rect 32456 44316 32462 44328
rect 32861 44319 32919 44325
rect 32861 44316 32873 44319
rect 32456 44288 32873 44316
rect 32456 44276 32462 44288
rect 32861 44285 32873 44288
rect 32907 44316 32919 44319
rect 32950 44316 32956 44328
rect 32907 44288 32956 44316
rect 32907 44285 32919 44288
rect 32861 44279 32919 44285
rect 32950 44276 32956 44288
rect 33008 44276 33014 44328
rect 33505 44319 33563 44325
rect 33505 44285 33517 44319
rect 33551 44285 33563 44319
rect 33505 44279 33563 44285
rect 31573 44251 31631 44257
rect 31573 44217 31585 44251
rect 31619 44248 31631 44251
rect 33520 44248 33548 44279
rect 34422 44276 34428 44328
rect 34480 44316 34486 44328
rect 35176 44316 35204 44347
rect 36630 44344 36636 44356
rect 36688 44344 36694 44396
rect 36909 44387 36967 44393
rect 36909 44353 36921 44387
rect 36955 44384 36967 44387
rect 37458 44384 37464 44396
rect 36955 44356 37464 44384
rect 36955 44353 36967 44356
rect 36909 44347 36967 44353
rect 37458 44344 37464 44356
rect 37516 44344 37522 44396
rect 38194 44384 38200 44396
rect 38155 44356 38200 44384
rect 38194 44344 38200 44356
rect 38252 44344 38258 44396
rect 38930 44384 38936 44396
rect 38891 44356 38936 44384
rect 38930 44344 38936 44356
rect 38988 44344 38994 44396
rect 39114 44384 39120 44396
rect 39075 44356 39120 44384
rect 39114 44344 39120 44356
rect 39172 44344 39178 44396
rect 40126 44344 40132 44396
rect 40184 44384 40190 44396
rect 40589 44387 40647 44393
rect 40589 44384 40601 44387
rect 40184 44356 40601 44384
rect 40184 44344 40190 44356
rect 40589 44353 40601 44356
rect 40635 44353 40647 44387
rect 42242 44384 42248 44396
rect 40589 44347 40647 44353
rect 40972 44356 42248 44384
rect 34480 44288 35204 44316
rect 36648 44316 36676 44344
rect 37182 44316 37188 44328
rect 36648 44288 37188 44316
rect 34480 44276 34486 44288
rect 37182 44276 37188 44288
rect 37240 44276 37246 44328
rect 37734 44276 37740 44328
rect 37792 44316 37798 44328
rect 37918 44316 37924 44328
rect 37792 44288 37924 44316
rect 37792 44276 37798 44288
rect 37918 44276 37924 44288
rect 37976 44276 37982 44328
rect 38102 44316 38108 44328
rect 38063 44288 38108 44316
rect 38102 44276 38108 44288
rect 38160 44276 38166 44328
rect 39945 44319 40003 44325
rect 39945 44285 39957 44319
rect 39991 44316 40003 44319
rect 40681 44319 40739 44325
rect 40681 44316 40693 44319
rect 39991 44288 40693 44316
rect 39991 44285 40003 44288
rect 39945 44279 40003 44285
rect 40681 44285 40693 44288
rect 40727 44316 40739 44319
rect 40862 44316 40868 44328
rect 40727 44288 40868 44316
rect 40727 44285 40739 44288
rect 40681 44279 40739 44285
rect 40862 44276 40868 44288
rect 40920 44276 40926 44328
rect 36906 44248 36912 44260
rect 31619 44220 33548 44248
rect 36867 44220 36912 44248
rect 31619 44217 31631 44220
rect 31573 44211 31631 44217
rect 36906 44208 36912 44220
rect 36964 44208 36970 44260
rect 40972 44248 41000 44356
rect 42242 44344 42248 44356
rect 42300 44344 42306 44396
rect 42426 44344 42432 44396
rect 42484 44384 42490 44396
rect 42613 44387 42671 44393
rect 42613 44384 42625 44387
rect 42484 44356 42625 44384
rect 42484 44344 42490 44356
rect 42613 44353 42625 44356
rect 42659 44353 42671 44387
rect 42886 44384 42892 44396
rect 42799 44356 42892 44384
rect 42613 44347 42671 44353
rect 42886 44344 42892 44356
rect 42944 44344 42950 44396
rect 43640 44393 43668 44424
rect 44450 44412 44456 44424
rect 44508 44412 44514 44464
rect 47210 44412 47216 44464
rect 47268 44452 47274 44464
rect 48148 44461 48176 44492
rect 48406 44480 48412 44492
rect 48464 44480 48470 44532
rect 48498 44480 48504 44532
rect 48556 44520 48562 44532
rect 49234 44520 49240 44532
rect 48556 44492 49240 44520
rect 48556 44480 48562 44492
rect 49234 44480 49240 44492
rect 49292 44480 49298 44532
rect 48133 44455 48191 44461
rect 47268 44424 47901 44452
rect 47268 44412 47274 44424
rect 43625 44387 43683 44393
rect 43625 44353 43637 44387
rect 43671 44353 43683 44387
rect 43625 44347 43683 44353
rect 46845 44387 46903 44393
rect 46845 44353 46857 44387
rect 46891 44384 46903 44387
rect 46934 44384 46940 44396
rect 46891 44356 46940 44384
rect 46891 44353 46903 44356
rect 46845 44347 46903 44353
rect 46934 44344 46940 44356
rect 46992 44344 46998 44396
rect 47121 44387 47179 44393
rect 47121 44353 47133 44387
rect 47167 44384 47179 44387
rect 47302 44384 47308 44396
rect 47167 44356 47308 44384
rect 47167 44353 47179 44356
rect 47121 44347 47179 44353
rect 47302 44344 47308 44356
rect 47360 44344 47366 44396
rect 47873 44393 47901 44424
rect 48133 44421 48145 44455
rect 48179 44452 48191 44455
rect 49145 44455 49203 44461
rect 48179 44424 49005 44452
rect 48179 44421 48191 44424
rect 48133 44415 48191 44421
rect 48977 44396 49005 44424
rect 49145 44421 49157 44455
rect 49191 44452 49203 44455
rect 51166 44452 51172 44464
rect 49191 44424 51172 44452
rect 49191 44421 49203 44424
rect 49145 44415 49203 44421
rect 47765 44387 47823 44393
rect 47765 44353 47777 44387
rect 47811 44353 47823 44387
rect 47765 44347 47823 44353
rect 47858 44387 47916 44393
rect 47858 44353 47870 44387
rect 47904 44353 47916 44387
rect 47858 44347 47916 44353
rect 48041 44387 48099 44393
rect 48041 44353 48053 44387
rect 48087 44384 48099 44387
rect 48271 44387 48329 44393
rect 48087 44356 48176 44384
rect 48087 44353 48099 44356
rect 48041 44347 48099 44353
rect 41506 44276 41512 44328
rect 41564 44316 41570 44328
rect 42904 44316 42932 44344
rect 43530 44316 43536 44328
rect 41564 44288 42932 44316
rect 43491 44288 43536 44316
rect 41564 44276 41570 44288
rect 43530 44276 43536 44288
rect 43588 44276 43594 44328
rect 43990 44316 43996 44328
rect 43951 44288 43996 44316
rect 43990 44276 43996 44288
rect 44048 44276 44054 44328
rect 37016 44220 41000 44248
rect 32214 44140 32220 44192
rect 32272 44180 32278 44192
rect 32582 44180 32588 44192
rect 32272 44152 32588 44180
rect 32272 44140 32278 44152
rect 32582 44140 32588 44152
rect 32640 44180 32646 44192
rect 32677 44183 32735 44189
rect 32677 44180 32689 44183
rect 32640 44152 32689 44180
rect 32640 44140 32646 44152
rect 32677 44149 32689 44152
rect 32723 44149 32735 44183
rect 32677 44143 32735 44149
rect 36722 44140 36728 44192
rect 36780 44180 36786 44192
rect 37016 44180 37044 44220
rect 41230 44208 41236 44260
rect 41288 44248 41294 44260
rect 41288 44220 42104 44248
rect 41288 44208 41294 44220
rect 38010 44180 38016 44192
rect 36780 44152 37044 44180
rect 37971 44152 38016 44180
rect 36780 44140 36786 44152
rect 38010 44140 38016 44152
rect 38068 44140 38074 44192
rect 38378 44140 38384 44192
rect 38436 44180 38442 44192
rect 39206 44180 39212 44192
rect 38436 44152 39212 44180
rect 38436 44140 38442 44152
rect 39206 44140 39212 44152
rect 39264 44140 39270 44192
rect 40678 44140 40684 44192
rect 40736 44180 40742 44192
rect 40957 44183 41015 44189
rect 40957 44180 40969 44183
rect 40736 44152 40969 44180
rect 40736 44140 40742 44152
rect 40957 44149 40969 44152
rect 41003 44149 41015 44183
rect 42076 44180 42104 44220
rect 42150 44208 42156 44260
rect 42208 44248 42214 44260
rect 42613 44251 42671 44257
rect 42613 44248 42625 44251
rect 42208 44220 42625 44248
rect 42208 44208 42214 44220
rect 42613 44217 42625 44220
rect 42659 44217 42671 44251
rect 42613 44211 42671 44217
rect 46845 44251 46903 44257
rect 46845 44217 46857 44251
rect 46891 44248 46903 44251
rect 47780 44248 47808 44347
rect 46891 44220 47808 44248
rect 46891 44217 46903 44220
rect 46845 44211 46903 44217
rect 48148 44192 48176 44356
rect 48271 44353 48283 44387
rect 48317 44353 48329 44387
rect 48866 44384 48872 44396
rect 48827 44356 48872 44384
rect 48271 44347 48329 44353
rect 48286 44316 48314 44347
rect 48866 44344 48872 44356
rect 48924 44344 48930 44396
rect 48958 44344 48964 44396
rect 49016 44384 49022 44396
rect 49234 44384 49240 44396
rect 49016 44356 49061 44384
rect 49195 44356 49240 44384
rect 49016 44344 49022 44356
rect 49234 44344 49240 44356
rect 49292 44344 49298 44396
rect 49334 44387 49392 44393
rect 49334 44353 49346 44387
rect 49380 44353 49392 44387
rect 49334 44347 49392 44353
rect 49349 44316 49377 44347
rect 48286 44288 49377 44316
rect 48976 44260 49004 44288
rect 48958 44208 48964 44260
rect 49016 44208 49022 44260
rect 49436 44248 49464 44424
rect 51166 44412 51172 44424
rect 51224 44452 51230 44464
rect 51224 44424 52040 44452
rect 51224 44412 51230 44424
rect 50249 44387 50307 44393
rect 50249 44353 50261 44387
rect 50295 44353 50307 44387
rect 50430 44384 50436 44396
rect 50391 44356 50436 44384
rect 50249 44347 50307 44353
rect 50264 44316 50292 44347
rect 50430 44344 50436 44356
rect 50488 44344 50494 44396
rect 50525 44387 50583 44393
rect 50525 44353 50537 44387
rect 50571 44384 50583 44387
rect 51718 44384 51724 44396
rect 50571 44356 51120 44384
rect 51679 44356 51724 44384
rect 50571 44353 50583 44356
rect 50525 44347 50583 44353
rect 50982 44316 50988 44328
rect 50264 44288 50988 44316
rect 50982 44276 50988 44288
rect 51040 44276 51046 44328
rect 51092 44316 51120 44356
rect 51718 44344 51724 44356
rect 51776 44344 51782 44396
rect 52012 44393 52040 44424
rect 52086 44412 52092 44464
rect 52144 44452 52150 44464
rect 52144 44424 52189 44452
rect 52144 44412 52150 44424
rect 51814 44387 51872 44393
rect 51814 44353 51826 44387
rect 51860 44353 51872 44387
rect 51814 44347 51872 44353
rect 51997 44387 52055 44393
rect 51997 44353 52009 44387
rect 52043 44353 52055 44387
rect 51997 44347 52055 44353
rect 52227 44387 52285 44393
rect 52227 44353 52239 44387
rect 52273 44384 52285 44387
rect 52822 44384 52828 44396
rect 52273 44356 52828 44384
rect 52273 44353 52285 44356
rect 52227 44347 52285 44353
rect 51626 44316 51632 44328
rect 51092 44288 51632 44316
rect 51626 44276 51632 44288
rect 51684 44276 51690 44328
rect 49068 44220 49464 44248
rect 46290 44180 46296 44192
rect 42076 44152 46296 44180
rect 40957 44143 41015 44149
rect 46290 44140 46296 44152
rect 46348 44140 46354 44192
rect 47210 44140 47216 44192
rect 47268 44180 47274 44192
rect 48130 44180 48136 44192
rect 47268 44152 48136 44180
rect 47268 44140 47274 44152
rect 48130 44140 48136 44152
rect 48188 44180 48194 44192
rect 49068 44180 49096 44220
rect 50798 44208 50804 44260
rect 50856 44248 50862 44260
rect 51828 44248 51856 44347
rect 52012 44316 52040 44347
rect 52822 44344 52828 44356
rect 52880 44344 52886 44396
rect 53006 44384 53012 44396
rect 52967 44356 53012 44384
rect 53006 44344 53012 44356
rect 53064 44344 53070 44396
rect 53193 44387 53251 44393
rect 53193 44353 53205 44387
rect 53239 44353 53251 44387
rect 54570 44384 54576 44396
rect 54531 44356 54576 44384
rect 53193 44347 53251 44353
rect 52012 44288 52316 44316
rect 52288 44260 52316 44288
rect 50856 44220 51856 44248
rect 50856 44208 50862 44220
rect 52270 44208 52276 44260
rect 52328 44208 52334 44260
rect 52365 44251 52423 44257
rect 52365 44217 52377 44251
rect 52411 44248 52423 44251
rect 53208 44248 53236 44347
rect 54570 44344 54576 44356
rect 54628 44344 54634 44396
rect 54941 44387 54999 44393
rect 54941 44353 54953 44387
rect 54987 44384 54999 44387
rect 55766 44384 55772 44396
rect 54987 44356 55772 44384
rect 54987 44353 54999 44356
rect 54941 44347 54999 44353
rect 54021 44319 54079 44325
rect 54021 44285 54033 44319
rect 54067 44316 54079 44319
rect 54956 44316 54984 44347
rect 55766 44344 55772 44356
rect 55824 44344 55830 44396
rect 54067 44288 54984 44316
rect 55585 44319 55643 44325
rect 54067 44285 54079 44288
rect 54021 44279 54079 44285
rect 55585 44285 55597 44319
rect 55631 44316 55643 44319
rect 56134 44316 56140 44328
rect 55631 44288 56140 44316
rect 55631 44285 55643 44288
rect 55585 44279 55643 44285
rect 56134 44276 56140 44288
rect 56192 44276 56198 44328
rect 52411 44220 53236 44248
rect 52411 44217 52423 44220
rect 52365 44211 52423 44217
rect 48188 44152 49096 44180
rect 48188 44140 48194 44152
rect 49234 44140 49240 44192
rect 49292 44180 49298 44192
rect 49513 44183 49571 44189
rect 49513 44180 49525 44183
rect 49292 44152 49525 44180
rect 49292 44140 49298 44152
rect 49513 44149 49525 44152
rect 49559 44149 49571 44183
rect 49513 44143 49571 44149
rect 50249 44183 50307 44189
rect 50249 44149 50261 44183
rect 50295 44180 50307 44183
rect 50338 44180 50344 44192
rect 50295 44152 50344 44180
rect 50295 44149 50307 44152
rect 50249 44143 50307 44149
rect 50338 44140 50344 44152
rect 50396 44140 50402 44192
rect 50522 44140 50528 44192
rect 50580 44180 50586 44192
rect 51077 44183 51135 44189
rect 51077 44180 51089 44183
rect 50580 44152 51089 44180
rect 50580 44140 50586 44152
rect 51077 44149 51089 44152
rect 51123 44180 51135 44183
rect 52638 44180 52644 44192
rect 51123 44152 52644 44180
rect 51123 44149 51135 44152
rect 51077 44143 51135 44149
rect 52638 44140 52644 44152
rect 52696 44140 52702 44192
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 34149 43979 34207 43985
rect 34149 43945 34161 43979
rect 34195 43976 34207 43979
rect 34238 43976 34244 43988
rect 34195 43948 34244 43976
rect 34195 43945 34207 43948
rect 34149 43939 34207 43945
rect 34238 43936 34244 43948
rect 34296 43936 34302 43988
rect 36354 43936 36360 43988
rect 36412 43976 36418 43988
rect 37090 43976 37096 43988
rect 36412 43948 37096 43976
rect 36412 43936 36418 43948
rect 37090 43936 37096 43948
rect 37148 43976 37154 43988
rect 41322 43976 41328 43988
rect 37148 43948 41328 43976
rect 37148 43936 37154 43948
rect 41322 43936 41328 43948
rect 41380 43976 41386 43988
rect 41509 43979 41567 43985
rect 41380 43936 41414 43976
rect 41509 43945 41521 43979
rect 41555 43976 41567 43979
rect 42702 43976 42708 43988
rect 41555 43948 42708 43976
rect 41555 43945 41567 43948
rect 41509 43939 41567 43945
rect 42702 43936 42708 43948
rect 42760 43936 42766 43988
rect 42797 43979 42855 43985
rect 42797 43945 42809 43979
rect 42843 43976 42855 43979
rect 43530 43976 43536 43988
rect 42843 43948 43536 43976
rect 42843 43945 42855 43948
rect 42797 43939 42855 43945
rect 43530 43936 43536 43948
rect 43588 43936 43594 43988
rect 43806 43936 43812 43988
rect 43864 43976 43870 43988
rect 46293 43979 46351 43985
rect 46293 43976 46305 43979
rect 43864 43948 46305 43976
rect 43864 43936 43870 43948
rect 46293 43945 46305 43948
rect 46339 43945 46351 43979
rect 46293 43939 46351 43945
rect 33318 43868 33324 43920
rect 33376 43908 33382 43920
rect 34885 43911 34943 43917
rect 34885 43908 34897 43911
rect 33376 43880 34897 43908
rect 33376 43868 33382 43880
rect 34885 43877 34897 43880
rect 34931 43908 34943 43911
rect 35342 43908 35348 43920
rect 34931 43880 35348 43908
rect 34931 43877 34943 43880
rect 34885 43871 34943 43877
rect 35342 43868 35348 43880
rect 35400 43908 35406 43920
rect 35529 43911 35587 43917
rect 35529 43908 35541 43911
rect 35400 43880 35541 43908
rect 35400 43868 35406 43880
rect 35529 43877 35541 43880
rect 35575 43877 35587 43911
rect 35529 43871 35587 43877
rect 36262 43868 36268 43920
rect 36320 43908 36326 43920
rect 36449 43911 36507 43917
rect 36449 43908 36461 43911
rect 36320 43880 36461 43908
rect 36320 43868 36326 43880
rect 36449 43877 36461 43880
rect 36495 43908 36507 43911
rect 41138 43908 41144 43920
rect 36495 43880 41144 43908
rect 36495 43877 36507 43880
rect 36449 43871 36507 43877
rect 41138 43868 41144 43880
rect 41196 43868 41202 43920
rect 41386 43908 41414 43936
rect 41386 43880 41920 43908
rect 32585 43843 32643 43849
rect 32585 43809 32597 43843
rect 32631 43840 32643 43843
rect 34422 43840 34428 43852
rect 32631 43812 34428 43840
rect 32631 43809 32643 43812
rect 32585 43803 32643 43809
rect 34422 43800 34428 43812
rect 34480 43800 34486 43852
rect 40678 43840 40684 43852
rect 37200 43812 38976 43840
rect 40639 43812 40684 43840
rect 31110 43732 31116 43784
rect 31168 43772 31174 43784
rect 31665 43775 31723 43781
rect 31665 43772 31677 43775
rect 31168 43744 31677 43772
rect 31168 43732 31174 43744
rect 31665 43741 31677 43744
rect 31711 43741 31723 43775
rect 31665 43735 31723 43741
rect 32033 43775 32091 43781
rect 32033 43741 32045 43775
rect 32079 43772 32091 43775
rect 32674 43772 32680 43784
rect 32079 43744 32680 43772
rect 32079 43741 32091 43744
rect 32033 43735 32091 43741
rect 32674 43732 32680 43744
rect 32732 43732 32738 43784
rect 37090 43772 37096 43784
rect 37051 43744 37096 43772
rect 37090 43732 37096 43744
rect 37148 43732 37154 43784
rect 33229 43707 33287 43713
rect 33229 43673 33241 43707
rect 33275 43704 33287 43707
rect 33594 43704 33600 43716
rect 33275 43676 33600 43704
rect 33275 43673 33287 43676
rect 33229 43667 33287 43673
rect 33594 43664 33600 43676
rect 33652 43704 33658 43716
rect 34330 43704 34336 43716
rect 33652 43676 34336 43704
rect 33652 43664 33658 43676
rect 34330 43664 34336 43676
rect 34388 43664 34394 43716
rect 35066 43664 35072 43716
rect 35124 43704 35130 43716
rect 36173 43707 36231 43713
rect 36173 43704 36185 43707
rect 35124 43676 36185 43704
rect 35124 43664 35130 43676
rect 36173 43673 36185 43676
rect 36219 43704 36231 43707
rect 37200 43704 37228 43812
rect 38010 43732 38016 43784
rect 38068 43772 38074 43784
rect 38289 43775 38347 43781
rect 38289 43772 38301 43775
rect 38068 43744 38301 43772
rect 38068 43732 38074 43744
rect 38289 43741 38301 43744
rect 38335 43741 38347 43775
rect 38289 43735 38347 43741
rect 38378 43732 38384 43784
rect 38436 43772 38442 43784
rect 38746 43772 38752 43784
rect 38804 43781 38810 43784
rect 38436 43744 38481 43772
rect 38712 43744 38752 43772
rect 38436 43732 38442 43744
rect 38746 43732 38752 43744
rect 38804 43735 38812 43781
rect 38948 43772 38976 43812
rect 40678 43800 40684 43812
rect 40736 43800 40742 43852
rect 41598 43840 41604 43852
rect 40788 43812 41604 43840
rect 40586 43772 40592 43784
rect 38948 43744 39988 43772
rect 40547 43744 40592 43772
rect 38804 43732 38810 43735
rect 36219 43676 37228 43704
rect 37461 43707 37519 43713
rect 36219 43673 36231 43676
rect 36173 43667 36231 43673
rect 37461 43673 37473 43707
rect 37507 43704 37519 43707
rect 38194 43704 38200 43716
rect 37507 43676 38200 43704
rect 37507 43673 37519 43676
rect 37461 43667 37519 43673
rect 38194 43664 38200 43676
rect 38252 43664 38258 43716
rect 38470 43664 38476 43716
rect 38528 43704 38534 43716
rect 38565 43707 38623 43713
rect 38565 43704 38577 43707
rect 38528 43676 38577 43704
rect 38528 43664 38534 43676
rect 38565 43673 38577 43676
rect 38611 43673 38623 43707
rect 38565 43667 38623 43673
rect 38657 43707 38715 43713
rect 38657 43673 38669 43707
rect 38703 43704 38715 43707
rect 39114 43704 39120 43716
rect 38703 43676 38884 43704
rect 38703 43673 38715 43676
rect 38657 43667 38715 43673
rect 38856 43648 38884 43676
rect 38948 43676 39120 43704
rect 33505 43639 33563 43645
rect 33505 43605 33517 43639
rect 33551 43636 33563 43639
rect 33778 43636 33784 43648
rect 33551 43608 33784 43636
rect 33551 43605 33563 43608
rect 33505 43599 33563 43605
rect 33778 43596 33784 43608
rect 33836 43636 33842 43648
rect 34054 43636 34060 43648
rect 33836 43608 34060 43636
rect 33836 43596 33842 43608
rect 34054 43596 34060 43608
rect 34112 43596 34118 43648
rect 38838 43596 38844 43648
rect 38896 43596 38902 43648
rect 38948 43645 38976 43676
rect 39114 43664 39120 43676
rect 39172 43664 39178 43716
rect 39960 43704 39988 43744
rect 40586 43732 40592 43744
rect 40644 43732 40650 43784
rect 40788 43704 40816 43812
rect 41598 43800 41604 43812
rect 41656 43800 41662 43852
rect 41693 43843 41751 43849
rect 41693 43809 41705 43843
rect 41739 43809 41751 43843
rect 41693 43803 41751 43809
rect 41417 43775 41475 43781
rect 41417 43741 41429 43775
rect 41463 43741 41475 43775
rect 41417 43735 41475 43741
rect 39960 43676 40816 43704
rect 41322 43664 41328 43716
rect 41380 43704 41386 43716
rect 41432 43704 41460 43735
rect 41506 43732 41512 43784
rect 41564 43772 41570 43784
rect 41708 43772 41736 43803
rect 41564 43744 41736 43772
rect 41564 43732 41570 43744
rect 41380 43676 41460 43704
rect 41892 43704 41920 43880
rect 42150 43868 42156 43920
rect 42208 43908 42214 43920
rect 45738 43908 45744 43920
rect 42208 43880 45600 43908
rect 45699 43880 45744 43908
rect 42208 43868 42214 43880
rect 42886 43840 42892 43852
rect 42444 43812 42892 43840
rect 41966 43732 41972 43784
rect 42024 43772 42030 43784
rect 42334 43781 42340 43784
rect 42153 43775 42211 43781
rect 42153 43772 42165 43775
rect 42024 43744 42165 43772
rect 42024 43732 42030 43744
rect 42153 43741 42165 43744
rect 42199 43741 42211 43775
rect 42153 43735 42211 43741
rect 42301 43775 42340 43781
rect 42301 43741 42313 43775
rect 42301 43735 42340 43741
rect 42334 43732 42340 43735
rect 42392 43732 42398 43784
rect 42444 43781 42472 43812
rect 42886 43800 42892 43812
rect 42944 43800 42950 43852
rect 45278 43840 45284 43852
rect 45239 43812 45284 43840
rect 45278 43800 45284 43812
rect 45336 43800 45342 43852
rect 45572 43840 45600 43880
rect 45738 43868 45744 43880
rect 45796 43868 45802 43920
rect 46308 43908 46336 43939
rect 46474 43936 46480 43988
rect 46532 43976 46538 43988
rect 46845 43979 46903 43985
rect 46845 43976 46857 43979
rect 46532 43948 46857 43976
rect 46532 43936 46538 43948
rect 46845 43945 46857 43948
rect 46891 43945 46903 43979
rect 50430 43976 50436 43988
rect 46845 43939 46903 43945
rect 47136 43948 50436 43976
rect 47026 43908 47032 43920
rect 46308 43880 47032 43908
rect 47026 43868 47032 43880
rect 47084 43868 47090 43920
rect 47136 43840 47164 43948
rect 50430 43936 50436 43948
rect 50488 43936 50494 43988
rect 50614 43936 50620 43988
rect 50672 43976 50678 43988
rect 50985 43979 51043 43985
rect 50985 43976 50997 43979
rect 50672 43948 50997 43976
rect 50672 43936 50678 43948
rect 50985 43945 50997 43948
rect 51031 43945 51043 43979
rect 50985 43939 51043 43945
rect 51629 43979 51687 43985
rect 51629 43945 51641 43979
rect 51675 43976 51687 43979
rect 51718 43976 51724 43988
rect 51675 43948 51724 43976
rect 51675 43945 51687 43948
rect 51629 43939 51687 43945
rect 51718 43936 51724 43948
rect 51776 43936 51782 43988
rect 54021 43979 54079 43985
rect 54021 43945 54033 43979
rect 54067 43976 54079 43979
rect 54570 43976 54576 43988
rect 54067 43948 54576 43976
rect 54067 43945 54079 43948
rect 54021 43939 54079 43945
rect 54570 43936 54576 43948
rect 54628 43936 54634 43988
rect 48222 43868 48228 43920
rect 48280 43908 48286 43920
rect 48280 43880 50752 43908
rect 48280 43868 48286 43880
rect 48958 43840 48964 43852
rect 45572 43812 47164 43840
rect 47320 43812 48964 43840
rect 42429 43775 42487 43781
rect 42429 43741 42441 43775
rect 42475 43741 42487 43775
rect 42429 43735 42487 43741
rect 42659 43775 42717 43781
rect 42659 43741 42671 43775
rect 42705 43772 42717 43775
rect 43070 43772 43076 43784
rect 42705 43744 43076 43772
rect 42705 43741 42717 43744
rect 42659 43735 42717 43741
rect 43070 43732 43076 43744
rect 43128 43772 43134 43784
rect 43257 43775 43315 43781
rect 43257 43772 43269 43775
rect 43128 43744 43269 43772
rect 43128 43732 43134 43744
rect 43257 43741 43269 43744
rect 43303 43741 43315 43775
rect 45370 43772 45376 43784
rect 45331 43744 45376 43772
rect 43257 43735 43315 43741
rect 45370 43732 45376 43744
rect 45428 43732 45434 43784
rect 47024 43775 47082 43781
rect 47024 43741 47036 43775
rect 47070 43772 47082 43775
rect 47320 43772 47348 43812
rect 48958 43800 48964 43812
rect 49016 43800 49022 43852
rect 49142 43840 49148 43852
rect 49103 43812 49148 43840
rect 49142 43800 49148 43812
rect 49200 43800 49206 43852
rect 49602 43800 49608 43852
rect 49660 43840 49666 43852
rect 50724 43840 50752 43880
rect 50798 43868 50804 43920
rect 50856 43908 50862 43920
rect 52457 43911 52515 43917
rect 52457 43908 52469 43911
rect 50856 43880 52469 43908
rect 50856 43868 50862 43880
rect 52457 43877 52469 43880
rect 52503 43908 52515 43911
rect 53926 43908 53932 43920
rect 52503 43880 53932 43908
rect 52503 43877 52515 43880
rect 52457 43871 52515 43877
rect 53926 43868 53932 43880
rect 53984 43868 53990 43920
rect 49660 43812 50660 43840
rect 50724 43812 51028 43840
rect 49660 43800 49666 43812
rect 47070 43744 47348 43772
rect 47396 43775 47454 43781
rect 47070 43741 47082 43744
rect 47024 43735 47082 43741
rect 47396 43741 47408 43775
rect 47442 43741 47454 43775
rect 47396 43735 47454 43741
rect 42518 43704 42524 43716
rect 41892 43676 42524 43704
rect 41380 43664 41386 43676
rect 42518 43664 42524 43676
rect 42576 43664 42582 43716
rect 44085 43707 44143 43713
rect 44085 43673 44097 43707
rect 44131 43704 44143 43707
rect 44266 43704 44272 43716
rect 44131 43676 44272 43704
rect 44131 43673 44143 43676
rect 44085 43667 44143 43673
rect 44266 43664 44272 43676
rect 44324 43664 44330 43716
rect 47118 43704 47124 43716
rect 47079 43676 47124 43704
rect 47118 43664 47124 43676
rect 47176 43664 47182 43716
rect 47210 43664 47216 43716
rect 47268 43704 47274 43716
rect 47412 43704 47440 43735
rect 47486 43732 47492 43784
rect 47544 43772 47550 43784
rect 49234 43772 49240 43784
rect 47544 43744 47589 43772
rect 49195 43744 49240 43772
rect 47544 43732 47550 43744
rect 49234 43732 49240 43744
rect 49292 43732 49298 43784
rect 50338 43772 50344 43784
rect 50299 43744 50344 43772
rect 50338 43732 50344 43744
rect 50396 43732 50402 43784
rect 50522 43781 50528 43784
rect 50489 43775 50528 43781
rect 50489 43741 50501 43775
rect 50489 43735 50528 43741
rect 50522 43732 50528 43735
rect 50580 43732 50586 43784
rect 50632 43772 50660 43812
rect 51000 43784 51028 43812
rect 51534 43800 51540 43852
rect 51592 43840 51598 43852
rect 53561 43843 53619 43849
rect 53561 43840 53573 43843
rect 51592 43812 53573 43840
rect 51592 43800 51598 43812
rect 53561 43809 53573 43812
rect 53607 43809 53619 43843
rect 53561 43803 53619 43809
rect 55490 43800 55496 43852
rect 55548 43840 55554 43852
rect 56505 43843 56563 43849
rect 56505 43840 56517 43843
rect 55548 43812 56517 43840
rect 55548 43800 55554 43812
rect 56505 43809 56517 43812
rect 56551 43809 56563 43843
rect 56505 43803 56563 43809
rect 50806 43775 50864 43781
rect 50806 43772 50818 43775
rect 50632 43744 50818 43772
rect 50806 43741 50818 43744
rect 50852 43741 50864 43775
rect 50806 43735 50864 43741
rect 50982 43732 50988 43784
rect 51040 43772 51046 43784
rect 51629 43775 51687 43781
rect 51629 43772 51641 43775
rect 51040 43744 51641 43772
rect 51040 43732 51046 43744
rect 51629 43741 51641 43744
rect 51675 43741 51687 43775
rect 51629 43735 51687 43741
rect 51810 43732 51816 43784
rect 51868 43772 51874 43784
rect 51905 43775 51963 43781
rect 51905 43772 51917 43775
rect 51868 43744 51917 43772
rect 51868 43732 51874 43744
rect 51905 43741 51917 43744
rect 51951 43741 51963 43775
rect 53650 43772 53656 43784
rect 53611 43744 53656 43772
rect 51905 43735 51963 43741
rect 53650 43732 53656 43744
rect 53708 43732 53714 43784
rect 55306 43732 55312 43784
rect 55364 43772 55370 43784
rect 55585 43775 55643 43781
rect 55585 43772 55597 43775
rect 55364 43744 55597 43772
rect 55364 43732 55370 43744
rect 55585 43741 55597 43744
rect 55631 43741 55643 43775
rect 55766 43772 55772 43784
rect 55727 43744 55772 43772
rect 55585 43735 55643 43741
rect 55766 43732 55772 43744
rect 55824 43732 55830 43784
rect 47670 43704 47676 43716
rect 47268 43676 47313 43704
rect 47412 43676 47676 43704
rect 47268 43664 47274 43676
rect 38933 43639 38991 43645
rect 38933 43605 38945 43639
rect 38979 43605 38991 43639
rect 38933 43599 38991 43605
rect 39022 43596 39028 43648
rect 39080 43636 39086 43648
rect 39390 43636 39396 43648
rect 39080 43608 39396 43636
rect 39080 43596 39086 43608
rect 39390 43596 39396 43608
rect 39448 43596 39454 43648
rect 40954 43636 40960 43648
rect 40915 43608 40960 43636
rect 40954 43596 40960 43608
rect 41012 43596 41018 43648
rect 41693 43639 41751 43645
rect 41693 43605 41705 43639
rect 41739 43636 41751 43639
rect 42610 43636 42616 43648
rect 41739 43608 42616 43636
rect 41739 43605 41751 43608
rect 41693 43599 41751 43605
rect 42610 43596 42616 43608
rect 42668 43596 42674 43648
rect 42978 43596 42984 43648
rect 43036 43636 43042 43648
rect 43441 43639 43499 43645
rect 43441 43636 43453 43639
rect 43036 43608 43453 43636
rect 43036 43596 43042 43608
rect 43441 43605 43453 43608
rect 43487 43636 43499 43639
rect 44174 43636 44180 43648
rect 43487 43608 44180 43636
rect 43487 43605 43499 43608
rect 43441 43599 43499 43605
rect 44174 43596 44180 43608
rect 44232 43596 44238 43648
rect 44542 43636 44548 43648
rect 44503 43608 44548 43636
rect 44542 43596 44548 43608
rect 44600 43596 44606 43648
rect 47026 43596 47032 43648
rect 47084 43636 47090 43648
rect 47412 43636 47440 43676
rect 47670 43664 47676 43676
rect 47728 43704 47734 43716
rect 48225 43707 48283 43713
rect 48225 43704 48237 43707
rect 47728 43676 48237 43704
rect 47728 43664 47734 43676
rect 48225 43673 48237 43676
rect 48271 43704 48283 43707
rect 48774 43704 48780 43716
rect 48271 43676 48780 43704
rect 48271 43673 48283 43676
rect 48225 43667 48283 43673
rect 48774 43664 48780 43676
rect 48832 43664 48838 43716
rect 50617 43707 50675 43713
rect 50617 43673 50629 43707
rect 50663 43673 50675 43707
rect 50617 43667 50675 43673
rect 48314 43636 48320 43648
rect 47084 43608 47440 43636
rect 48275 43608 48320 43636
rect 47084 43596 47090 43608
rect 48314 43596 48320 43608
rect 48372 43596 48378 43648
rect 49605 43639 49663 43645
rect 49605 43605 49617 43639
rect 49651 43636 49663 43639
rect 50062 43636 50068 43648
rect 49651 43608 50068 43636
rect 49651 43605 49663 43608
rect 49605 43599 49663 43605
rect 50062 43596 50068 43608
rect 50120 43596 50126 43648
rect 50632 43636 50660 43667
rect 50706 43664 50712 43716
rect 50764 43704 50770 43716
rect 55030 43704 55036 43716
rect 50764 43676 50809 43704
rect 52932 43676 55036 43704
rect 50764 43664 50770 43676
rect 50890 43636 50896 43648
rect 50632 43608 50896 43636
rect 50890 43596 50896 43608
rect 50948 43596 50954 43648
rect 51813 43639 51871 43645
rect 51813 43605 51825 43639
rect 51859 43636 51871 43639
rect 52086 43636 52092 43648
rect 51859 43608 52092 43636
rect 51859 43605 51871 43608
rect 51813 43599 51871 43605
rect 52086 43596 52092 43608
rect 52144 43636 52150 43648
rect 52932 43645 52960 43676
rect 55030 43664 55036 43676
rect 55088 43664 55094 43716
rect 52917 43639 52975 43645
rect 52917 43636 52929 43639
rect 52144 43608 52929 43636
rect 52144 43596 52150 43608
rect 52917 43605 52929 43608
rect 52963 43605 52975 43639
rect 52917 43599 52975 43605
rect 53282 43596 53288 43648
rect 53340 43636 53346 43648
rect 54478 43636 54484 43648
rect 53340 43608 54484 43636
rect 53340 43596 53346 43608
rect 54478 43596 54484 43608
rect 54536 43596 54542 43648
rect 1104 43546 58880 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 35594 43546
rect 35646 43494 35658 43546
rect 35710 43494 35722 43546
rect 35774 43494 35786 43546
rect 35838 43494 35850 43546
rect 35902 43494 58880 43546
rect 1104 43472 58880 43494
rect 34333 43435 34391 43441
rect 34333 43401 34345 43435
rect 34379 43432 34391 43435
rect 34514 43432 34520 43444
rect 34379 43404 34520 43432
rect 34379 43401 34391 43404
rect 34333 43395 34391 43401
rect 34514 43392 34520 43404
rect 34572 43392 34578 43444
rect 35342 43392 35348 43444
rect 35400 43432 35406 43444
rect 36078 43432 36084 43444
rect 35400 43404 36084 43432
rect 35400 43392 35406 43404
rect 36078 43392 36084 43404
rect 36136 43392 36142 43444
rect 36265 43435 36323 43441
rect 36265 43401 36277 43435
rect 36311 43432 36323 43435
rect 38565 43435 38623 43441
rect 36311 43404 37780 43432
rect 36311 43401 36323 43404
rect 36265 43395 36323 43401
rect 30745 43299 30803 43305
rect 30745 43265 30757 43299
rect 30791 43296 30803 43299
rect 31018 43296 31024 43308
rect 30791 43268 31024 43296
rect 30791 43265 30803 43268
rect 30745 43259 30803 43265
rect 31018 43256 31024 43268
rect 31076 43256 31082 43308
rect 32950 43296 32956 43308
rect 32911 43268 32956 43296
rect 32950 43256 32956 43268
rect 33008 43296 33014 43308
rect 33008 43268 33916 43296
rect 33008 43256 33014 43268
rect 30006 43188 30012 43240
rect 30064 43228 30070 43240
rect 30653 43231 30711 43237
rect 30653 43228 30665 43231
rect 30064 43200 30665 43228
rect 30064 43188 30070 43200
rect 30653 43197 30665 43200
rect 30699 43197 30711 43231
rect 31110 43228 31116 43240
rect 31071 43200 31116 43228
rect 30653 43191 30711 43197
rect 31110 43188 31116 43200
rect 31168 43188 31174 43240
rect 32858 43228 32864 43240
rect 32819 43200 32864 43228
rect 32858 43188 32864 43200
rect 32916 43188 32922 43240
rect 33888 43237 33916 43268
rect 33962 43256 33968 43308
rect 34020 43296 34026 43308
rect 34020 43268 34065 43296
rect 34020 43256 34026 43268
rect 34790 43256 34796 43308
rect 34848 43296 34854 43308
rect 34977 43299 35035 43305
rect 34977 43296 34989 43299
rect 34848 43268 34989 43296
rect 34848 43256 34854 43268
rect 34977 43265 34989 43268
rect 35023 43265 35035 43299
rect 34977 43259 35035 43265
rect 35066 43256 35072 43308
rect 35124 43296 35130 43308
rect 35250 43296 35256 43308
rect 35124 43268 35169 43296
rect 35211 43268 35256 43296
rect 35124 43256 35130 43268
rect 35250 43256 35256 43268
rect 35308 43256 35314 43308
rect 35365 43305 35393 43392
rect 36170 43324 36176 43376
rect 36228 43364 36234 43376
rect 36541 43367 36599 43373
rect 36541 43364 36553 43367
rect 36228 43336 36553 43364
rect 36228 43324 36234 43336
rect 36541 43333 36553 43336
rect 36587 43333 36599 43367
rect 36541 43327 36599 43333
rect 35526 43305 35532 43308
rect 35345 43299 35403 43305
rect 35345 43265 35357 43299
rect 35391 43265 35403 43299
rect 35345 43259 35403 43265
rect 35481 43299 35532 43305
rect 35481 43265 35493 43299
rect 35527 43265 35532 43299
rect 35481 43259 35532 43265
rect 35526 43256 35532 43259
rect 35584 43296 35590 43308
rect 36403 43299 36461 43305
rect 36403 43296 36415 43299
rect 35584 43268 36415 43296
rect 35584 43256 35590 43268
rect 36403 43265 36415 43268
rect 36449 43265 36461 43299
rect 36630 43296 36636 43308
rect 36591 43268 36636 43296
rect 36403 43259 36461 43265
rect 36630 43256 36636 43268
rect 36688 43256 36694 43308
rect 36722 43256 36728 43308
rect 36780 43305 36786 43308
rect 36780 43299 36819 43305
rect 36807 43265 36819 43299
rect 36780 43259 36819 43265
rect 36780 43256 36786 43259
rect 36906 43256 36912 43308
rect 36964 43296 36970 43308
rect 37752 43305 37780 43404
rect 38565 43401 38577 43435
rect 38611 43432 38623 43435
rect 40402 43432 40408 43444
rect 38611 43404 40408 43432
rect 38611 43401 38623 43404
rect 38565 43395 38623 43401
rect 40402 43392 40408 43404
rect 40460 43392 40466 43444
rect 40586 43432 40592 43444
rect 40547 43404 40592 43432
rect 40586 43392 40592 43404
rect 40644 43392 40650 43444
rect 41598 43392 41604 43444
rect 41656 43432 41662 43444
rect 41785 43435 41843 43441
rect 41785 43432 41797 43435
rect 41656 43404 41797 43432
rect 41656 43392 41662 43404
rect 41785 43401 41797 43404
rect 41831 43432 41843 43435
rect 42334 43432 42340 43444
rect 41831 43404 42340 43432
rect 41831 43401 41843 43404
rect 41785 43395 41843 43401
rect 42334 43392 42340 43404
rect 42392 43392 42398 43444
rect 42702 43432 42708 43444
rect 42444 43404 42708 43432
rect 39298 43364 39304 43376
rect 37844 43336 39304 43364
rect 37737 43299 37795 43305
rect 36964 43268 37009 43296
rect 36964 43256 36970 43268
rect 37737 43265 37749 43299
rect 37783 43265 37795 43299
rect 37737 43259 37795 43265
rect 33873 43231 33931 43237
rect 33873 43197 33885 43231
rect 33919 43197 33931 43231
rect 33873 43191 33931 43197
rect 34054 43188 34060 43240
rect 34112 43228 34118 43240
rect 35084 43228 35112 43256
rect 35618 43228 35624 43240
rect 34112 43200 35624 43228
rect 34112 43188 34118 43200
rect 35618 43188 35624 43200
rect 35676 43188 35682 43240
rect 37645 43231 37703 43237
rect 37645 43197 37657 43231
rect 37691 43197 37703 43231
rect 37645 43191 37703 43197
rect 33321 43163 33379 43169
rect 33321 43129 33333 43163
rect 33367 43160 33379 43163
rect 37660 43160 37688 43191
rect 33367 43132 37688 43160
rect 33367 43129 33379 43132
rect 33321 43123 33379 43129
rect 33962 43052 33968 43104
rect 34020 43092 34026 43104
rect 35621 43095 35679 43101
rect 35621 43092 35633 43095
rect 34020 43064 35633 43092
rect 34020 43052 34026 43064
rect 35621 43061 35633 43064
rect 35667 43061 35679 43095
rect 35621 43055 35679 43061
rect 36722 43052 36728 43104
rect 36780 43092 36786 43104
rect 37090 43092 37096 43104
rect 36780 43064 37096 43092
rect 36780 43052 36786 43064
rect 37090 43052 37096 43064
rect 37148 43092 37154 43104
rect 37844 43092 37872 43336
rect 39298 43324 39304 43336
rect 39356 43324 39362 43376
rect 39485 43367 39543 43373
rect 39485 43333 39497 43367
rect 39531 43333 39543 43367
rect 39485 43327 39543 43333
rect 41972 43367 42030 43373
rect 41972 43333 41984 43367
rect 42018 43364 42030 43367
rect 42444 43364 42472 43404
rect 42702 43392 42708 43404
rect 42760 43392 42766 43444
rect 43257 43435 43315 43441
rect 43257 43401 43269 43435
rect 43303 43432 43315 43435
rect 43438 43432 43444 43444
rect 43303 43404 43444 43432
rect 43303 43401 43315 43404
rect 43257 43395 43315 43401
rect 43438 43392 43444 43404
rect 43496 43392 43502 43444
rect 44361 43435 44419 43441
rect 44361 43401 44373 43435
rect 44407 43401 44419 43435
rect 46290 43432 46296 43444
rect 46251 43404 46296 43432
rect 44361 43395 44419 43401
rect 42018 43336 42472 43364
rect 42018 43333 42030 43336
rect 41972 43327 42030 43333
rect 39206 43256 39212 43308
rect 39264 43296 39270 43308
rect 39500 43296 39528 43327
rect 42518 43324 42524 43376
rect 42576 43364 42582 43376
rect 42886 43364 42892 43376
rect 42576 43336 42749 43364
rect 42847 43336 42892 43364
rect 42576 43324 42582 43336
rect 39945 43299 40003 43305
rect 39945 43296 39957 43299
rect 39264 43268 39309 43296
rect 39500 43268 39957 43296
rect 39264 43256 39270 43268
rect 39945 43265 39957 43268
rect 39991 43265 40003 43299
rect 39945 43259 40003 43265
rect 40034 43256 40040 43308
rect 40092 43296 40098 43308
rect 40218 43296 40224 43308
rect 40092 43268 40137 43296
rect 40179 43268 40224 43296
rect 40092 43256 40098 43268
rect 40218 43256 40224 43268
rect 40276 43256 40282 43308
rect 40310 43256 40316 43308
rect 40368 43296 40374 43308
rect 40451 43299 40509 43305
rect 40368 43268 40413 43296
rect 40368 43256 40374 43268
rect 40451 43265 40463 43299
rect 40497 43296 40509 43299
rect 40678 43296 40684 43308
rect 40497 43268 40684 43296
rect 40497 43265 40509 43268
rect 40451 43259 40509 43265
rect 40678 43256 40684 43268
rect 40736 43256 40742 43308
rect 41690 43296 41696 43308
rect 41651 43268 41696 43296
rect 41690 43256 41696 43268
rect 41748 43256 41754 43308
rect 41782 43256 41788 43308
rect 41840 43296 41846 43308
rect 42610 43296 42616 43308
rect 41840 43268 42473 43296
rect 42571 43268 42616 43296
rect 41840 43256 41846 43268
rect 39482 43228 39488 43240
rect 39443 43200 39488 43228
rect 39482 43188 39488 43200
rect 39540 43228 39546 43240
rect 39758 43228 39764 43240
rect 39540 43200 39764 43228
rect 39540 43188 39546 43200
rect 39758 43188 39764 43200
rect 39816 43188 39822 43240
rect 41800 43228 41828 43256
rect 41156 43200 41828 43228
rect 42445 43228 42473 43268
rect 42610 43256 42616 43268
rect 42668 43256 42674 43308
rect 42721 43305 42749 43336
rect 42886 43324 42892 43336
rect 42944 43324 42950 43376
rect 43622 43324 43628 43376
rect 43680 43364 43686 43376
rect 43993 43367 44051 43373
rect 43993 43364 44005 43367
rect 43680 43336 44005 43364
rect 43680 43324 43686 43336
rect 43993 43333 44005 43336
rect 44039 43333 44051 43367
rect 43993 43327 44051 43333
rect 44085 43367 44143 43373
rect 44085 43333 44097 43367
rect 44131 43364 44143 43367
rect 44266 43364 44272 43376
rect 44131 43336 44272 43364
rect 44131 43333 44143 43336
rect 44085 43327 44143 43333
rect 44266 43324 44272 43336
rect 44324 43324 44330 43376
rect 42706 43299 42764 43305
rect 42706 43265 42718 43299
rect 42752 43265 42764 43299
rect 42706 43259 42764 43265
rect 42981 43299 43039 43305
rect 42981 43265 42993 43299
rect 43027 43265 43039 43299
rect 42981 43259 43039 43265
rect 42996 43228 43024 43259
rect 43070 43256 43076 43308
rect 43128 43305 43134 43308
rect 43128 43296 43136 43305
rect 43714 43296 43720 43308
rect 43128 43268 43173 43296
rect 43675 43268 43720 43296
rect 43128 43259 43136 43268
rect 43128 43256 43134 43259
rect 43714 43256 43720 43268
rect 43772 43256 43778 43308
rect 43898 43305 43904 43308
rect 43865 43299 43904 43305
rect 43865 43265 43877 43299
rect 43865 43259 43904 43265
rect 43898 43256 43904 43259
rect 43956 43256 43962 43308
rect 44174 43256 44180 43308
rect 44232 43305 44238 43308
rect 44232 43296 44240 43305
rect 44376 43296 44404 43395
rect 46290 43392 46296 43404
rect 46348 43392 46354 43444
rect 47121 43435 47179 43441
rect 47121 43401 47133 43435
rect 47167 43432 47179 43435
rect 47486 43432 47492 43444
rect 47167 43404 47492 43432
rect 47167 43401 47179 43404
rect 47121 43395 47179 43401
rect 47486 43392 47492 43404
rect 47544 43392 47550 43444
rect 47946 43392 47952 43444
rect 48004 43432 48010 43444
rect 48133 43435 48191 43441
rect 48133 43432 48145 43435
rect 48004 43404 48145 43432
rect 48004 43392 48010 43404
rect 48133 43401 48145 43404
rect 48179 43432 48191 43435
rect 48498 43432 48504 43444
rect 48179 43404 48504 43432
rect 48179 43401 48191 43404
rect 48133 43395 48191 43401
rect 48498 43392 48504 43404
rect 48556 43392 48562 43444
rect 52086 43432 52092 43444
rect 51046 43404 52092 43432
rect 51046 43364 51074 43404
rect 52086 43392 52092 43404
rect 52144 43392 52150 43444
rect 53926 43392 53932 43444
rect 53984 43432 53990 43444
rect 54021 43435 54079 43441
rect 54021 43432 54033 43435
rect 53984 43404 54033 43432
rect 53984 43392 53990 43404
rect 54021 43401 54033 43404
rect 54067 43432 54079 43435
rect 54294 43432 54300 43444
rect 54067 43404 54300 43432
rect 54067 43401 54079 43404
rect 54021 43395 54079 43401
rect 54294 43392 54300 43404
rect 54352 43392 54358 43444
rect 45112 43336 51074 43364
rect 45005 43299 45063 43305
rect 45005 43296 45017 43299
rect 44232 43268 44277 43296
rect 44376 43268 45017 43296
rect 44232 43259 44240 43268
rect 45005 43265 45017 43268
rect 45051 43265 45063 43299
rect 45005 43259 45063 43265
rect 44232 43256 44238 43259
rect 42445 43200 43024 43228
rect 38194 43120 38200 43172
rect 38252 43160 38258 43172
rect 41046 43160 41052 43172
rect 38252 43132 39436 43160
rect 38252 43120 38258 43132
rect 39298 43092 39304 43104
rect 37148 43064 37872 43092
rect 39259 43064 39304 43092
rect 37148 43052 37154 43064
rect 39298 43052 39304 43064
rect 39356 43052 39362 43104
rect 39408 43092 39436 43132
rect 40236 43132 41052 43160
rect 40236 43092 40264 43132
rect 41046 43120 41052 43132
rect 41104 43120 41110 43172
rect 39408 43064 40264 43092
rect 40310 43052 40316 43104
rect 40368 43092 40374 43104
rect 41156 43101 41184 43200
rect 44358 43188 44364 43240
rect 44416 43228 44422 43240
rect 44913 43231 44971 43237
rect 44913 43228 44925 43231
rect 44416 43200 44925 43228
rect 44416 43188 44422 43200
rect 44913 43197 44925 43200
rect 44959 43197 44971 43231
rect 44913 43191 44971 43197
rect 41966 43120 41972 43172
rect 42024 43160 42030 43172
rect 42024 43132 42069 43160
rect 42024 43120 42030 43132
rect 43714 43120 43720 43172
rect 43772 43160 43778 43172
rect 44174 43160 44180 43172
rect 43772 43132 44180 43160
rect 43772 43120 43778 43132
rect 44174 43120 44180 43132
rect 44232 43120 44238 43172
rect 41141 43095 41199 43101
rect 41141 43092 41153 43095
rect 40368 43064 41153 43092
rect 40368 43052 40374 43064
rect 41141 43061 41153 43064
rect 41187 43061 41199 43095
rect 41141 43055 41199 43061
rect 41506 43052 41512 43104
rect 41564 43092 41570 43104
rect 45112 43092 45140 43336
rect 46845 43299 46903 43305
rect 46845 43265 46857 43299
rect 46891 43296 46903 43299
rect 47026 43296 47032 43308
rect 46891 43268 47032 43296
rect 46891 43265 46903 43268
rect 46845 43259 46903 43265
rect 47026 43256 47032 43268
rect 47084 43256 47090 43308
rect 47302 43296 47308 43308
rect 47136 43268 47308 43296
rect 47136 43237 47164 43268
rect 47302 43256 47308 43268
rect 47360 43296 47366 43308
rect 48041 43299 48099 43305
rect 48041 43296 48053 43299
rect 47360 43268 48053 43296
rect 47360 43256 47366 43268
rect 48041 43265 48053 43268
rect 48087 43265 48099 43299
rect 48041 43259 48099 43265
rect 48222 43256 48228 43308
rect 48280 43296 48286 43308
rect 48317 43299 48375 43305
rect 48317 43296 48329 43299
rect 48280 43268 48329 43296
rect 48280 43256 48286 43268
rect 48317 43265 48329 43268
rect 48363 43265 48375 43299
rect 48317 43259 48375 43265
rect 48590 43256 48596 43308
rect 48648 43296 48654 43308
rect 48777 43299 48835 43305
rect 48777 43296 48789 43299
rect 48648 43268 48789 43296
rect 48648 43256 48654 43268
rect 48777 43265 48789 43268
rect 48823 43296 48835 43299
rect 49602 43296 49608 43308
rect 48823 43268 49608 43296
rect 48823 43265 48835 43268
rect 48777 43259 48835 43265
rect 49602 43256 49608 43268
rect 49660 43256 49666 43308
rect 50062 43296 50068 43308
rect 49975 43268 50068 43296
rect 50062 43256 50068 43268
rect 50120 43296 50126 43308
rect 50522 43296 50528 43308
rect 50120 43268 50528 43296
rect 50120 43256 50126 43268
rect 50522 43256 50528 43268
rect 50580 43256 50586 43308
rect 51534 43296 51540 43308
rect 51495 43268 51540 43296
rect 51534 43256 51540 43268
rect 51592 43256 51598 43308
rect 54938 43296 54944 43308
rect 54899 43268 54944 43296
rect 54938 43256 54944 43268
rect 54996 43256 55002 43308
rect 47121 43231 47179 43237
rect 47121 43197 47133 43231
rect 47167 43197 47179 43231
rect 49970 43228 49976 43240
rect 49931 43200 49976 43228
rect 47121 43191 47179 43197
rect 49970 43188 49976 43200
rect 50028 43188 50034 43240
rect 51261 43231 51319 43237
rect 51261 43228 51273 43231
rect 51046 43200 51273 43228
rect 45370 43160 45376 43172
rect 45331 43132 45376 43160
rect 45370 43120 45376 43132
rect 45428 43120 45434 43172
rect 46290 43120 46296 43172
rect 46348 43160 46354 43172
rect 47946 43160 47952 43172
rect 46348 43132 47952 43160
rect 46348 43120 46354 43132
rect 47946 43120 47952 43132
rect 48004 43120 48010 43172
rect 48317 43163 48375 43169
rect 48317 43129 48329 43163
rect 48363 43160 48375 43163
rect 48866 43160 48872 43172
rect 48363 43132 48872 43160
rect 48363 43129 48375 43132
rect 48317 43123 48375 43129
rect 48866 43120 48872 43132
rect 48924 43120 48930 43172
rect 50433 43163 50491 43169
rect 50433 43129 50445 43163
rect 50479 43160 50491 43163
rect 51046 43160 51074 43200
rect 51261 43197 51273 43200
rect 51307 43197 51319 43231
rect 51261 43191 51319 43197
rect 51442 43188 51448 43240
rect 51500 43228 51506 43240
rect 52089 43231 52147 43237
rect 52089 43228 52101 43231
rect 51500 43200 52101 43228
rect 51500 43188 51506 43200
rect 52089 43197 52101 43200
rect 52135 43197 52147 43231
rect 52089 43191 52147 43197
rect 55033 43231 55091 43237
rect 55033 43197 55045 43231
rect 55079 43197 55091 43231
rect 55306 43228 55312 43240
rect 55267 43200 55312 43228
rect 55033 43191 55091 43197
rect 52822 43160 52828 43172
rect 50479 43132 51074 43160
rect 51276 43132 52828 43160
rect 50479 43129 50491 43132
rect 50433 43123 50491 43129
rect 46934 43092 46940 43104
rect 41564 43064 45140 43092
rect 46847 43064 46940 43092
rect 41564 43052 41570 43064
rect 46934 43052 46940 43064
rect 46992 43092 46998 43104
rect 48222 43092 48228 43104
rect 46992 43064 48228 43092
rect 46992 43052 46998 43064
rect 48222 43052 48228 43064
rect 48280 43052 48286 43104
rect 48958 43092 48964 43104
rect 48871 43064 48964 43092
rect 48958 43052 48964 43064
rect 49016 43092 49022 43104
rect 51276 43092 51304 43132
rect 52822 43120 52828 43132
rect 52880 43120 52886 43172
rect 55048 43160 55076 43191
rect 55306 43188 55312 43200
rect 55364 43188 55370 43240
rect 55214 43160 55220 43172
rect 55048 43132 55220 43160
rect 55214 43120 55220 43132
rect 55272 43120 55278 43172
rect 49016 43064 51304 43092
rect 49016 43052 49022 43064
rect 52638 43052 52644 43104
rect 52696 43092 52702 43104
rect 52917 43095 52975 43101
rect 52917 43092 52929 43095
rect 52696 43064 52929 43092
rect 52696 43052 52702 43064
rect 52917 43061 52929 43064
rect 52963 43092 52975 43095
rect 53466 43092 53472 43104
rect 52963 43064 53472 43092
rect 52963 43061 52975 43064
rect 52917 43055 52975 43061
rect 53466 43052 53472 43064
rect 53524 43052 53530 43104
rect 55122 43052 55128 43104
rect 55180 43092 55186 43104
rect 55769 43095 55827 43101
rect 55769 43092 55781 43095
rect 55180 43064 55781 43092
rect 55180 43052 55186 43064
rect 55769 43061 55781 43064
rect 55815 43061 55827 43095
rect 55769 43055 55827 43061
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 31113 42891 31171 42897
rect 31113 42857 31125 42891
rect 31159 42888 31171 42891
rect 32950 42888 32956 42900
rect 31159 42860 32956 42888
rect 31159 42857 31171 42860
rect 31113 42851 31171 42857
rect 32950 42848 32956 42860
rect 33008 42848 33014 42900
rect 33229 42891 33287 42897
rect 33229 42857 33241 42891
rect 33275 42888 33287 42891
rect 33318 42888 33324 42900
rect 33275 42860 33324 42888
rect 33275 42857 33287 42860
rect 33229 42851 33287 42857
rect 32674 42820 32680 42832
rect 32635 42792 32680 42820
rect 32674 42780 32680 42792
rect 32732 42780 32738 42832
rect 30190 42712 30196 42764
rect 30248 42752 30254 42764
rect 30745 42755 30803 42761
rect 30745 42752 30757 42755
rect 30248 42724 30757 42752
rect 30248 42712 30254 42724
rect 30745 42721 30757 42724
rect 30791 42721 30803 42755
rect 30745 42715 30803 42721
rect 31846 42712 31852 42764
rect 31904 42752 31910 42764
rect 33244 42752 33272 42851
rect 33318 42848 33324 42860
rect 33376 42848 33382 42900
rect 36446 42888 36452 42900
rect 35177 42860 36452 42888
rect 34149 42823 34207 42829
rect 34149 42789 34161 42823
rect 34195 42820 34207 42823
rect 34698 42820 34704 42832
rect 34195 42792 34704 42820
rect 34195 42789 34207 42792
rect 34149 42783 34207 42789
rect 34698 42780 34704 42792
rect 34756 42780 34762 42832
rect 31904 42724 32168 42752
rect 31904 42712 31910 42724
rect 30837 42687 30895 42693
rect 30837 42653 30849 42687
rect 30883 42684 30895 42687
rect 31386 42684 31392 42696
rect 30883 42656 31392 42684
rect 30883 42653 30895 42656
rect 30837 42647 30895 42653
rect 31386 42644 31392 42656
rect 31444 42644 31450 42696
rect 31754 42644 31760 42696
rect 31812 42684 31818 42696
rect 32140 42693 32168 42724
rect 32416 42724 33272 42752
rect 34333 42755 34391 42761
rect 32033 42687 32091 42693
rect 32033 42684 32045 42687
rect 31812 42656 32045 42684
rect 31812 42644 31818 42656
rect 32033 42653 32045 42656
rect 32079 42653 32091 42687
rect 32033 42647 32091 42653
rect 32126 42687 32184 42693
rect 32126 42653 32138 42687
rect 32172 42684 32184 42687
rect 32214 42684 32220 42696
rect 32172 42656 32220 42684
rect 32172 42653 32184 42656
rect 32126 42647 32184 42653
rect 32214 42644 32220 42656
rect 32272 42644 32278 42696
rect 32416 42693 32444 42724
rect 34333 42721 34345 42755
rect 34379 42752 34391 42755
rect 34974 42752 34980 42764
rect 34379 42724 34980 42752
rect 34379 42721 34391 42724
rect 34333 42715 34391 42721
rect 34974 42712 34980 42724
rect 35032 42712 35038 42764
rect 32401 42687 32459 42693
rect 32401 42653 32413 42687
rect 32447 42653 32459 42687
rect 32401 42647 32459 42653
rect 32490 42644 32496 42696
rect 32548 42693 32554 42696
rect 32548 42684 32556 42693
rect 34054 42684 34060 42696
rect 32548 42656 32593 42684
rect 34015 42656 34060 42684
rect 32548 42647 32556 42656
rect 32548 42644 32554 42647
rect 34054 42644 34060 42656
rect 34112 42644 34118 42696
rect 35177 42693 35205 42860
rect 36446 42848 36452 42860
rect 36504 42848 36510 42900
rect 36906 42848 36912 42900
rect 36964 42888 36970 42900
rect 37001 42891 37059 42897
rect 37001 42888 37013 42891
rect 36964 42860 37013 42888
rect 36964 42848 36970 42860
rect 37001 42857 37013 42860
rect 37047 42857 37059 42891
rect 37001 42851 37059 42857
rect 37090 42848 37096 42900
rect 37148 42888 37154 42900
rect 40218 42888 40224 42900
rect 37148 42860 37193 42888
rect 37292 42860 40224 42888
rect 37148 42848 37154 42860
rect 36357 42823 36415 42829
rect 36357 42789 36369 42823
rect 36403 42789 36415 42823
rect 36357 42783 36415 42789
rect 36372 42752 36400 42783
rect 36630 42780 36636 42832
rect 36688 42820 36694 42832
rect 37292 42820 37320 42860
rect 40218 42848 40224 42860
rect 40276 42888 40282 42900
rect 40402 42888 40408 42900
rect 40276 42860 40408 42888
rect 40276 42848 40282 42860
rect 40402 42848 40408 42860
rect 40460 42848 40466 42900
rect 41966 42848 41972 42900
rect 42024 42888 42030 42900
rect 42794 42888 42800 42900
rect 42024 42860 42800 42888
rect 42024 42848 42030 42860
rect 42794 42848 42800 42860
rect 42852 42888 42858 42900
rect 42889 42891 42947 42897
rect 42889 42888 42901 42891
rect 42852 42860 42901 42888
rect 42852 42848 42858 42860
rect 42889 42857 42901 42860
rect 42935 42888 42947 42891
rect 43438 42888 43444 42900
rect 42935 42860 43444 42888
rect 42935 42857 42947 42860
rect 42889 42851 42947 42857
rect 43438 42848 43444 42860
rect 43496 42888 43502 42900
rect 44361 42891 44419 42897
rect 44361 42888 44373 42891
rect 43496 42860 44373 42888
rect 43496 42848 43502 42860
rect 44361 42857 44373 42860
rect 44407 42857 44419 42891
rect 47210 42888 47216 42900
rect 44361 42851 44419 42857
rect 46400 42860 47216 42888
rect 36688 42792 37320 42820
rect 38565 42823 38623 42829
rect 36688 42780 36694 42792
rect 38565 42789 38577 42823
rect 38611 42820 38623 42823
rect 38838 42820 38844 42832
rect 38611 42792 38844 42820
rect 38611 42789 38623 42792
rect 38565 42783 38623 42789
rect 38838 42780 38844 42792
rect 38896 42780 38902 42832
rect 39390 42780 39396 42832
rect 39448 42820 39454 42832
rect 43806 42820 43812 42832
rect 39448 42792 43812 42820
rect 39448 42780 39454 42792
rect 43806 42780 43812 42792
rect 43864 42780 43870 42832
rect 44634 42780 44640 42832
rect 44692 42820 44698 42832
rect 46400 42820 46428 42860
rect 47210 42848 47216 42860
rect 47268 42888 47274 42900
rect 48314 42888 48320 42900
rect 47268 42860 48320 42888
rect 47268 42848 47274 42860
rect 48314 42848 48320 42860
rect 48372 42848 48378 42900
rect 48406 42848 48412 42900
rect 48464 42888 48470 42900
rect 48501 42891 48559 42897
rect 48501 42888 48513 42891
rect 48464 42860 48513 42888
rect 48464 42848 48470 42860
rect 48501 42857 48513 42860
rect 48547 42857 48559 42891
rect 48501 42851 48559 42857
rect 48593 42891 48651 42897
rect 48593 42857 48605 42891
rect 48639 42888 48651 42891
rect 48866 42888 48872 42900
rect 48639 42860 48872 42888
rect 48639 42857 48651 42860
rect 48593 42851 48651 42857
rect 48866 42848 48872 42860
rect 48924 42848 48930 42900
rect 49789 42891 49847 42897
rect 49789 42857 49801 42891
rect 49835 42888 49847 42891
rect 49970 42888 49976 42900
rect 49835 42860 49976 42888
rect 49835 42857 49847 42860
rect 49789 42851 49847 42857
rect 49970 42848 49976 42860
rect 50028 42848 50034 42900
rect 53650 42848 53656 42900
rect 53708 42888 53714 42900
rect 53745 42891 53803 42897
rect 53745 42888 53757 42891
rect 53708 42860 53757 42888
rect 53708 42848 53714 42860
rect 53745 42857 53757 42860
rect 53791 42857 53803 42891
rect 53745 42851 53803 42857
rect 54849 42891 54907 42897
rect 54849 42857 54861 42891
rect 54895 42888 54907 42891
rect 54938 42888 54944 42900
rect 54895 42860 54944 42888
rect 54895 42857 54907 42860
rect 54849 42851 54907 42857
rect 54938 42848 54944 42860
rect 54996 42848 55002 42900
rect 44692 42792 46428 42820
rect 44692 42780 44698 42792
rect 47118 42780 47124 42832
rect 47176 42820 47182 42832
rect 49602 42820 49608 42832
rect 47176 42792 49608 42820
rect 47176 42780 47182 42792
rect 36909 42755 36967 42761
rect 36909 42752 36921 42755
rect 36372 42724 36921 42752
rect 36909 42721 36921 42724
rect 36955 42752 36967 42755
rect 37090 42752 37096 42764
rect 36955 42724 37096 42752
rect 36955 42721 36967 42724
rect 36909 42715 36967 42721
rect 37090 42712 37096 42724
rect 37148 42712 37154 42764
rect 37918 42712 37924 42764
rect 37976 42752 37982 42764
rect 38105 42755 38163 42761
rect 38105 42752 38117 42755
rect 37976 42724 38117 42752
rect 37976 42712 37982 42724
rect 38105 42721 38117 42724
rect 38151 42721 38163 42755
rect 38105 42715 38163 42721
rect 39298 42712 39304 42764
rect 39356 42752 39362 42764
rect 39666 42752 39672 42764
rect 39356 42724 39672 42752
rect 39356 42712 39362 42724
rect 39666 42712 39672 42724
rect 39724 42712 39730 42764
rect 44177 42755 44235 42761
rect 44177 42752 44189 42755
rect 42168 42724 44189 42752
rect 35069 42687 35127 42693
rect 35069 42653 35081 42687
rect 35115 42653 35127 42687
rect 35069 42647 35127 42653
rect 35162 42687 35220 42693
rect 35162 42653 35174 42687
rect 35208 42653 35220 42687
rect 35162 42647 35220 42653
rect 32309 42619 32367 42625
rect 32309 42585 32321 42619
rect 32355 42616 32367 42619
rect 33042 42616 33048 42628
rect 32355 42588 33048 42616
rect 32355 42585 32367 42588
rect 32309 42579 32367 42585
rect 33042 42576 33048 42588
rect 33100 42576 33106 42628
rect 34333 42619 34391 42625
rect 34333 42585 34345 42619
rect 34379 42616 34391 42619
rect 35084 42616 35112 42647
rect 35250 42644 35256 42696
rect 35308 42684 35314 42696
rect 35526 42684 35532 42696
rect 35584 42693 35590 42696
rect 35308 42656 35532 42684
rect 35308 42644 35314 42656
rect 35526 42644 35532 42656
rect 35584 42647 35592 42693
rect 35584 42644 35590 42647
rect 35986 42644 35992 42696
rect 36044 42684 36050 42696
rect 36173 42687 36231 42693
rect 36173 42684 36185 42687
rect 36044 42656 36185 42684
rect 36044 42644 36050 42656
rect 36173 42653 36185 42656
rect 36219 42653 36231 42687
rect 36173 42647 36231 42653
rect 37185 42687 37243 42693
rect 37185 42653 37197 42687
rect 37231 42653 37243 42687
rect 37185 42647 37243 42653
rect 35342 42616 35348 42628
rect 34379 42588 35112 42616
rect 35255 42588 35348 42616
rect 34379 42585 34391 42588
rect 34333 42579 34391 42585
rect 35342 42576 35348 42588
rect 35400 42576 35406 42628
rect 35437 42619 35495 42625
rect 35437 42585 35449 42619
rect 35483 42616 35495 42619
rect 35618 42616 35624 42628
rect 35483 42588 35624 42616
rect 35483 42585 35495 42588
rect 35437 42579 35495 42585
rect 35618 42576 35624 42588
rect 35676 42576 35682 42628
rect 34882 42508 34888 42560
rect 34940 42548 34946 42560
rect 35360 42548 35388 42576
rect 37200 42560 37228 42647
rect 37826 42644 37832 42696
rect 37884 42684 37890 42696
rect 38197 42687 38255 42693
rect 38197 42684 38209 42687
rect 37884 42656 38209 42684
rect 37884 42644 37890 42656
rect 38197 42653 38209 42656
rect 38243 42653 38255 42687
rect 38197 42647 38255 42653
rect 41782 42644 41788 42696
rect 41840 42684 41846 42696
rect 41969 42687 42027 42693
rect 41969 42684 41981 42687
rect 41840 42656 41981 42684
rect 41840 42644 41846 42656
rect 41969 42653 41981 42656
rect 42015 42653 42027 42687
rect 41969 42647 42027 42653
rect 34940 42520 35388 42548
rect 34940 42508 34946 42520
rect 35526 42508 35532 42560
rect 35584 42548 35590 42560
rect 35713 42551 35771 42557
rect 35713 42548 35725 42551
rect 35584 42520 35725 42548
rect 35584 42508 35590 42520
rect 35713 42517 35725 42520
rect 35759 42517 35771 42551
rect 35713 42511 35771 42517
rect 36170 42508 36176 42560
rect 36228 42548 36234 42560
rect 37182 42548 37188 42560
rect 36228 42520 37188 42548
rect 36228 42508 36234 42520
rect 37182 42508 37188 42520
rect 37240 42508 37246 42560
rect 38010 42508 38016 42560
rect 38068 42548 38074 42560
rect 38378 42548 38384 42560
rect 38068 42520 38384 42548
rect 38068 42508 38074 42520
rect 38378 42508 38384 42520
rect 38436 42548 38442 42560
rect 39025 42551 39083 42557
rect 39025 42548 39037 42551
rect 38436 42520 39037 42548
rect 38436 42508 38442 42520
rect 39025 42517 39037 42520
rect 39071 42517 39083 42551
rect 40034 42548 40040 42560
rect 39995 42520 40040 42548
rect 39025 42511 39083 42517
rect 40034 42508 40040 42520
rect 40092 42508 40098 42560
rect 41690 42508 41696 42560
rect 41748 42548 41754 42560
rect 42168 42557 42196 42724
rect 42702 42684 42708 42696
rect 42663 42656 42708 42684
rect 42702 42644 42708 42656
rect 42760 42644 42766 42696
rect 43438 42684 43444 42696
rect 43399 42656 43444 42684
rect 43438 42644 43444 42656
rect 43496 42644 43502 42696
rect 43732 42693 43760 42724
rect 44177 42721 44189 42724
rect 44223 42721 44235 42755
rect 44177 42715 44235 42721
rect 44266 42712 44272 42764
rect 44324 42752 44330 42764
rect 45002 42752 45008 42764
rect 44324 42724 45008 42752
rect 44324 42712 44330 42724
rect 45002 42712 45008 42724
rect 45060 42752 45066 42764
rect 48682 42752 48688 42764
rect 45060 42724 47716 42752
rect 48643 42724 48688 42752
rect 45060 42712 45066 42724
rect 43717 42687 43775 42693
rect 43717 42653 43729 42687
rect 43763 42653 43775 42687
rect 43717 42647 43775 42653
rect 43898 42644 43904 42696
rect 43956 42684 43962 42696
rect 44358 42684 44364 42696
rect 43956 42656 44364 42684
rect 43956 42644 43962 42656
rect 44358 42644 44364 42656
rect 44416 42684 44422 42696
rect 44453 42687 44511 42693
rect 44453 42684 44465 42687
rect 44416 42656 44465 42684
rect 44416 42644 44422 42656
rect 44453 42653 44465 42656
rect 44499 42684 44511 42687
rect 44542 42684 44548 42696
rect 44499 42656 44548 42684
rect 44499 42653 44511 42656
rect 44453 42647 44511 42653
rect 44542 42644 44548 42656
rect 44600 42644 44606 42696
rect 45554 42644 45560 42696
rect 45612 42684 45618 42696
rect 45741 42687 45799 42693
rect 45741 42684 45753 42687
rect 45612 42656 45753 42684
rect 45612 42644 45618 42656
rect 45741 42653 45753 42656
rect 45787 42653 45799 42687
rect 45741 42647 45799 42653
rect 45925 42687 45983 42693
rect 45925 42653 45937 42687
rect 45971 42653 45983 42687
rect 45925 42647 45983 42653
rect 44174 42616 44180 42628
rect 44135 42588 44180 42616
rect 44174 42576 44180 42588
rect 44232 42576 44238 42628
rect 44266 42576 44272 42628
rect 44324 42616 44330 42628
rect 45940 42616 45968 42647
rect 47688 42625 47716 42724
rect 48682 42712 48688 42724
rect 48740 42712 48746 42764
rect 48038 42644 48044 42696
rect 48096 42684 48102 42696
rect 48409 42687 48467 42693
rect 48409 42684 48421 42687
rect 48096 42656 48421 42684
rect 48096 42644 48102 42656
rect 48409 42653 48421 42656
rect 48455 42653 48467 42687
rect 48409 42647 48467 42653
rect 44324 42588 45968 42616
rect 46753 42619 46811 42625
rect 44324 42576 44330 42588
rect 46753 42585 46765 42619
rect 46799 42585 46811 42619
rect 46753 42579 46811 42585
rect 47673 42619 47731 42625
rect 47673 42585 47685 42619
rect 47719 42616 47731 42619
rect 48222 42616 48228 42628
rect 47719 42588 48228 42616
rect 47719 42585 47731 42588
rect 47673 42579 47731 42585
rect 42153 42551 42211 42557
rect 42153 42548 42165 42551
rect 41748 42520 42165 42548
rect 41748 42508 41754 42520
rect 42153 42517 42165 42520
rect 42199 42517 42211 42551
rect 42153 42511 42211 42517
rect 43346 42508 43352 42560
rect 43404 42548 43410 42560
rect 43539 42551 43597 42557
rect 43539 42548 43551 42551
rect 43404 42520 43551 42548
rect 43404 42508 43410 42520
rect 43539 42517 43551 42520
rect 43585 42517 43597 42551
rect 43539 42511 43597 42517
rect 43625 42551 43683 42557
rect 43625 42517 43637 42551
rect 43671 42548 43683 42551
rect 43714 42548 43720 42560
rect 43671 42520 43720 42548
rect 43671 42517 43683 42520
rect 43625 42511 43683 42517
rect 43714 42508 43720 42520
rect 43772 42508 43778 42560
rect 46768 42548 46796 42579
rect 48222 42576 48228 42588
rect 48280 42576 48286 42628
rect 48424 42616 48452 42647
rect 48866 42644 48872 42696
rect 48924 42684 48930 42696
rect 49253 42693 49281 42792
rect 49602 42780 49608 42792
rect 49660 42780 49666 42832
rect 52365 42823 52423 42829
rect 52365 42789 52377 42823
rect 52411 42820 52423 42823
rect 55214 42820 55220 42832
rect 52411 42792 55220 42820
rect 52411 42789 52423 42792
rect 52365 42783 52423 42789
rect 55214 42780 55220 42792
rect 55272 42820 55278 42832
rect 56413 42823 56471 42829
rect 55272 42792 56088 42820
rect 55272 42780 55278 42792
rect 51258 42712 51264 42764
rect 51316 42752 51322 42764
rect 51905 42755 51963 42761
rect 51905 42752 51917 42755
rect 51316 42724 51917 42752
rect 51316 42712 51322 42724
rect 51905 42721 51917 42724
rect 51951 42721 51963 42755
rect 51905 42715 51963 42721
rect 53374 42712 53380 42764
rect 53432 42752 53438 42764
rect 53432 42724 54248 42752
rect 53432 42712 53438 42724
rect 49145 42687 49203 42693
rect 49145 42684 49157 42687
rect 48924 42656 49157 42684
rect 48924 42644 48930 42656
rect 49145 42653 49157 42656
rect 49191 42653 49203 42687
rect 49145 42647 49203 42653
rect 49238 42687 49296 42693
rect 49238 42653 49250 42687
rect 49284 42653 49296 42687
rect 49418 42684 49424 42696
rect 49379 42656 49424 42684
rect 49238 42647 49296 42653
rect 49418 42644 49424 42656
rect 49476 42644 49482 42696
rect 49651 42687 49709 42693
rect 49651 42653 49663 42687
rect 49697 42684 49709 42687
rect 49878 42684 49884 42696
rect 49697 42656 49884 42684
rect 49697 42653 49709 42656
rect 49651 42647 49709 42653
rect 49878 42644 49884 42656
rect 49936 42644 49942 42696
rect 51994 42684 52000 42696
rect 51955 42656 52000 42684
rect 51994 42644 52000 42656
rect 52052 42644 52058 42696
rect 53098 42684 53104 42696
rect 53059 42656 53104 42684
rect 53098 42644 53104 42656
rect 53156 42644 53162 42696
rect 53194 42687 53252 42693
rect 53194 42653 53206 42687
rect 53240 42684 53252 42687
rect 53282 42684 53288 42696
rect 53240 42656 53288 42684
rect 53240 42653 53252 42656
rect 53194 42647 53252 42653
rect 49326 42616 49332 42628
rect 48424 42588 49332 42616
rect 49326 42576 49332 42588
rect 49384 42616 49390 42628
rect 49513 42619 49571 42625
rect 49513 42616 49525 42619
rect 49384 42588 49525 42616
rect 49384 42576 49390 42588
rect 49513 42585 49525 42588
rect 49559 42585 49571 42619
rect 50338 42616 50344 42628
rect 50299 42588 50344 42616
rect 49513 42579 49571 42585
rect 50338 42576 50344 42588
rect 50396 42616 50402 42628
rect 50893 42619 50951 42625
rect 50893 42616 50905 42619
rect 50396 42588 50905 42616
rect 50396 42576 50402 42588
rect 50893 42585 50905 42588
rect 50939 42616 50951 42619
rect 53208 42616 53236 42647
rect 53282 42644 53288 42656
rect 53340 42644 53346 42696
rect 53466 42684 53472 42696
rect 53427 42656 53472 42684
rect 53466 42644 53472 42656
rect 53524 42644 53530 42696
rect 53650 42693 53656 42696
rect 53607 42687 53656 42693
rect 53607 42653 53619 42687
rect 53653 42653 53656 42687
rect 53607 42647 53656 42653
rect 53650 42644 53656 42647
rect 53708 42644 53714 42696
rect 54220 42693 54248 42724
rect 54294 42712 54300 42764
rect 54352 42752 54358 42764
rect 54352 42724 54616 42752
rect 54352 42712 54358 42724
rect 54205 42687 54263 42693
rect 54205 42653 54217 42687
rect 54251 42653 54263 42687
rect 54386 42684 54392 42696
rect 54347 42656 54392 42684
rect 54205 42647 54263 42653
rect 54386 42644 54392 42656
rect 54444 42644 54450 42696
rect 54588 42693 54616 42724
rect 54754 42712 54760 42764
rect 54812 42752 54818 42764
rect 55953 42755 56011 42761
rect 55953 42752 55965 42755
rect 54812 42724 55965 42752
rect 54812 42712 54818 42724
rect 55953 42721 55965 42724
rect 55999 42721 56011 42755
rect 55953 42715 56011 42721
rect 54481 42687 54539 42693
rect 54481 42653 54493 42687
rect 54527 42653 54539 42687
rect 54481 42647 54539 42653
rect 54573 42687 54631 42693
rect 54573 42653 54585 42687
rect 54619 42684 54631 42687
rect 55122 42684 55128 42696
rect 54619 42656 55128 42684
rect 54619 42653 54631 42656
rect 54573 42647 54631 42653
rect 50939 42588 53236 42616
rect 53377 42619 53435 42625
rect 50939 42585 50951 42588
rect 50893 42579 50951 42585
rect 53377 42585 53389 42619
rect 53423 42585 53435 42619
rect 53377 42579 53435 42585
rect 49234 42548 49240 42560
rect 46768 42520 49240 42548
rect 49234 42508 49240 42520
rect 49292 42508 49298 42560
rect 51718 42508 51724 42560
rect 51776 42548 51782 42560
rect 53392 42548 53420 42579
rect 53742 42576 53748 42628
rect 53800 42616 53806 42628
rect 54496 42616 54524 42647
rect 55122 42644 55128 42656
rect 55180 42644 55186 42696
rect 56060 42693 56088 42792
rect 56413 42789 56425 42823
rect 56459 42820 56471 42823
rect 56459 42792 57192 42820
rect 56459 42789 56471 42792
rect 56413 42783 56471 42789
rect 57164 42761 57192 42792
rect 57149 42755 57207 42761
rect 57149 42721 57161 42755
rect 57195 42721 57207 42755
rect 57149 42715 57207 42721
rect 56045 42687 56103 42693
rect 56045 42653 56057 42687
rect 56091 42653 56103 42687
rect 57238 42684 57244 42696
rect 57199 42656 57244 42684
rect 56045 42647 56103 42653
rect 57238 42644 57244 42656
rect 57296 42644 57302 42696
rect 53800 42588 54524 42616
rect 53800 42576 53806 42588
rect 53926 42548 53932 42560
rect 51776 42520 53932 42548
rect 51776 42508 51782 42520
rect 53926 42508 53932 42520
rect 53984 42508 53990 42560
rect 54478 42508 54484 42560
rect 54536 42548 54542 42560
rect 56686 42548 56692 42560
rect 54536 42520 56692 42548
rect 54536 42508 54542 42520
rect 56686 42508 56692 42520
rect 56744 42508 56750 42560
rect 57054 42508 57060 42560
rect 57112 42548 57118 42560
rect 58069 42551 58127 42557
rect 58069 42548 58081 42551
rect 57112 42520 58081 42548
rect 57112 42508 57118 42520
rect 58069 42517 58081 42520
rect 58115 42517 58127 42551
rect 58069 42511 58127 42517
rect 1104 42458 58880 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 35594 42458
rect 35646 42406 35658 42458
rect 35710 42406 35722 42458
rect 35774 42406 35786 42458
rect 35838 42406 35850 42458
rect 35902 42406 58880 42458
rect 1104 42384 58880 42406
rect 31754 42304 31760 42356
rect 31812 42344 31818 42356
rect 31812 42316 31857 42344
rect 31812 42304 31818 42316
rect 32214 42304 32220 42356
rect 32272 42344 32278 42356
rect 32493 42347 32551 42353
rect 32493 42344 32505 42347
rect 32272 42316 32505 42344
rect 32272 42304 32278 42316
rect 32493 42313 32505 42316
rect 32539 42313 32551 42347
rect 32493 42307 32551 42313
rect 32508 42276 32536 42307
rect 34790 42304 34796 42356
rect 34848 42344 34854 42356
rect 34885 42347 34943 42353
rect 34885 42344 34897 42347
rect 34848 42316 34897 42344
rect 34848 42304 34854 42316
rect 34885 42313 34897 42316
rect 34931 42313 34943 42347
rect 34885 42307 34943 42313
rect 34974 42304 34980 42356
rect 35032 42344 35038 42356
rect 35986 42344 35992 42356
rect 35032 42316 35992 42344
rect 35032 42304 35038 42316
rect 35986 42304 35992 42316
rect 36044 42304 36050 42356
rect 36446 42304 36452 42356
rect 36504 42344 36510 42356
rect 36541 42347 36599 42353
rect 36541 42344 36553 42347
rect 36504 42316 36553 42344
rect 36504 42304 36510 42316
rect 36541 42313 36553 42316
rect 36587 42344 36599 42347
rect 36587 42316 37964 42344
rect 36587 42313 36599 42316
rect 36541 42307 36599 42313
rect 36170 42276 36176 42288
rect 32508 42248 36176 42276
rect 36170 42236 36176 42248
rect 36228 42236 36234 42288
rect 37936 42276 37964 42316
rect 38010 42304 38016 42356
rect 38068 42344 38074 42356
rect 39761 42347 39819 42353
rect 39761 42344 39773 42347
rect 38068 42316 39773 42344
rect 38068 42304 38074 42316
rect 39761 42313 39773 42316
rect 39807 42313 39819 42347
rect 43993 42347 44051 42353
rect 39761 42307 39819 42313
rect 42812 42316 43760 42344
rect 37936 42248 41460 42276
rect 29825 42211 29883 42217
rect 29825 42177 29837 42211
rect 29871 42208 29883 42211
rect 30006 42208 30012 42220
rect 29871 42180 30012 42208
rect 29871 42177 29883 42180
rect 29825 42171 29883 42177
rect 30006 42168 30012 42180
rect 30064 42168 30070 42220
rect 31110 42168 31116 42220
rect 31168 42208 31174 42220
rect 31481 42211 31539 42217
rect 31481 42208 31493 42211
rect 31168 42180 31493 42208
rect 31168 42168 31174 42180
rect 31481 42177 31493 42180
rect 31527 42208 31539 42211
rect 32214 42208 32220 42220
rect 31527 42180 32220 42208
rect 31527 42177 31539 42180
rect 31481 42171 31539 42177
rect 32214 42168 32220 42180
rect 32272 42208 32278 42220
rect 32401 42211 32459 42217
rect 32401 42208 32413 42211
rect 32272 42180 32413 42208
rect 32272 42168 32278 42180
rect 32401 42177 32413 42180
rect 32447 42177 32459 42211
rect 32401 42171 32459 42177
rect 34146 42168 34152 42220
rect 34204 42208 34210 42220
rect 34606 42208 34612 42220
rect 34204 42180 34612 42208
rect 34204 42168 34210 42180
rect 34606 42168 34612 42180
rect 34664 42168 34670 42220
rect 34698 42168 34704 42220
rect 34756 42208 34762 42220
rect 35713 42211 35771 42217
rect 34756 42180 34801 42208
rect 34756 42168 34762 42180
rect 35713 42177 35725 42211
rect 35759 42208 35771 42211
rect 36078 42208 36084 42220
rect 35759 42180 36084 42208
rect 35759 42177 35771 42180
rect 35713 42171 35771 42177
rect 36078 42168 36084 42180
rect 36136 42208 36142 42220
rect 36265 42211 36323 42217
rect 36265 42208 36277 42211
rect 36136 42180 36277 42208
rect 36136 42168 36142 42180
rect 36265 42177 36277 42180
rect 36311 42177 36323 42211
rect 36265 42171 36323 42177
rect 37461 42211 37519 42217
rect 37461 42177 37473 42211
rect 37507 42177 37519 42211
rect 38930 42208 38936 42220
rect 38891 42180 38936 42208
rect 37461 42171 37519 42177
rect 29270 42100 29276 42152
rect 29328 42140 29334 42152
rect 29733 42143 29791 42149
rect 29733 42140 29745 42143
rect 29328 42112 29745 42140
rect 29328 42100 29334 42112
rect 29733 42109 29745 42112
rect 29779 42109 29791 42143
rect 30190 42140 30196 42152
rect 30151 42112 30196 42140
rect 29733 42103 29791 42109
rect 30190 42100 30196 42112
rect 30248 42100 30254 42152
rect 31757 42143 31815 42149
rect 31757 42109 31769 42143
rect 31803 42140 31815 42143
rect 34885 42143 34943 42149
rect 31803 42112 32444 42140
rect 31803 42109 31815 42112
rect 31757 42103 31815 42109
rect 32416 42084 32444 42112
rect 34885 42109 34897 42143
rect 34931 42140 34943 42143
rect 34974 42140 34980 42152
rect 34931 42112 34980 42140
rect 34931 42109 34943 42112
rect 34885 42103 34943 42109
rect 34974 42100 34980 42112
rect 35032 42140 35038 42152
rect 35342 42140 35348 42152
rect 35032 42112 35348 42140
rect 35032 42100 35038 42112
rect 35342 42100 35348 42112
rect 35400 42100 35406 42152
rect 35434 42100 35440 42152
rect 35492 42140 35498 42152
rect 37476 42140 37504 42171
rect 38930 42168 38936 42180
rect 38988 42168 38994 42220
rect 40589 42211 40647 42217
rect 40589 42177 40601 42211
rect 40635 42208 40647 42211
rect 40770 42208 40776 42220
rect 40635 42180 40776 42208
rect 40635 42177 40647 42180
rect 40589 42171 40647 42177
rect 40770 42168 40776 42180
rect 40828 42168 40834 42220
rect 38838 42140 38844 42152
rect 35492 42112 37504 42140
rect 38799 42112 38844 42140
rect 35492 42100 35498 42112
rect 38838 42100 38844 42112
rect 38896 42100 38902 42152
rect 40497 42143 40555 42149
rect 40497 42140 40509 42143
rect 38948 42112 40509 42140
rect 32398 42032 32404 42084
rect 32456 42032 32462 42084
rect 33686 42032 33692 42084
rect 33744 42072 33750 42084
rect 38948 42072 38976 42112
rect 40497 42109 40509 42112
rect 40543 42109 40555 42143
rect 41432 42140 41460 42248
rect 41506 42236 41512 42288
rect 41564 42276 41570 42288
rect 42061 42279 42119 42285
rect 42061 42276 42073 42279
rect 41564 42248 42073 42276
rect 41564 42236 41570 42248
rect 42061 42245 42073 42248
rect 42107 42276 42119 42279
rect 42702 42276 42708 42288
rect 42107 42248 42708 42276
rect 42107 42245 42119 42248
rect 42061 42239 42119 42245
rect 42702 42236 42708 42248
rect 42760 42236 42766 42288
rect 41782 42208 41788 42220
rect 41743 42180 41788 42208
rect 41782 42168 41788 42180
rect 41840 42168 41846 42220
rect 41874 42168 41880 42220
rect 41932 42208 41938 42220
rect 41932 42180 41977 42208
rect 41932 42168 41938 42180
rect 42812 42149 42840 42316
rect 43732 42285 43760 42316
rect 43993 42313 44005 42347
rect 44039 42344 44051 42347
rect 44266 42344 44272 42356
rect 44039 42316 44272 42344
rect 44039 42313 44051 42316
rect 43993 42307 44051 42313
rect 44266 42304 44272 42316
rect 44324 42304 44330 42356
rect 45554 42344 45560 42356
rect 45515 42316 45560 42344
rect 45554 42304 45560 42316
rect 45612 42304 45618 42356
rect 47121 42347 47179 42353
rect 47121 42313 47133 42347
rect 47167 42344 47179 42347
rect 47210 42344 47216 42356
rect 47167 42316 47216 42344
rect 47167 42313 47179 42316
rect 47121 42307 47179 42313
rect 47210 42304 47216 42316
rect 47268 42304 47274 42356
rect 48958 42344 48964 42356
rect 47959 42316 48964 42344
rect 43717 42279 43775 42285
rect 43717 42245 43729 42279
rect 43763 42276 43775 42279
rect 47854 42276 47860 42288
rect 43763 42248 47860 42276
rect 43763 42245 43775 42248
rect 43717 42239 43775 42245
rect 47854 42236 47860 42248
rect 47912 42236 47918 42288
rect 43346 42208 43352 42220
rect 43307 42180 43352 42208
rect 43346 42168 43352 42180
rect 43404 42168 43410 42220
rect 43442 42211 43500 42217
rect 43442 42177 43454 42211
rect 43488 42208 43500 42211
rect 43530 42208 43536 42220
rect 43488 42180 43536 42208
rect 43488 42177 43500 42180
rect 43442 42171 43500 42177
rect 43530 42168 43536 42180
rect 43588 42168 43594 42220
rect 43622 42168 43628 42220
rect 43680 42208 43686 42220
rect 43898 42217 43904 42220
rect 43855 42211 43904 42217
rect 43680 42180 43773 42208
rect 43680 42168 43686 42180
rect 43855 42177 43867 42211
rect 43901 42177 43904 42211
rect 43855 42171 43904 42177
rect 43898 42168 43904 42171
rect 43956 42168 43962 42220
rect 45189 42211 45247 42217
rect 45189 42208 45201 42211
rect 44008 42180 45201 42208
rect 42797 42143 42855 42149
rect 42797 42140 42809 42143
rect 41432 42112 42809 42140
rect 40497 42103 40555 42109
rect 42797 42109 42809 42112
rect 42843 42109 42855 42143
rect 42797 42103 42855 42109
rect 42978 42100 42984 42152
rect 43036 42140 43042 42152
rect 43640 42140 43668 42168
rect 43036 42112 43668 42140
rect 43036 42100 43042 42112
rect 39298 42072 39304 42084
rect 33744 42044 38976 42072
rect 39259 42044 39304 42072
rect 33744 42032 33750 42044
rect 39298 42032 39304 42044
rect 39356 42032 39362 42084
rect 40957 42075 41015 42081
rect 40957 42041 40969 42075
rect 41003 42072 41015 42075
rect 41003 42044 42472 42072
rect 41003 42041 41015 42044
rect 40957 42035 41015 42041
rect 31573 42007 31631 42013
rect 31573 41973 31585 42007
rect 31619 42004 31631 42007
rect 32674 42004 32680 42016
rect 31619 41976 32680 42004
rect 31619 41973 31631 41976
rect 31573 41967 31631 41973
rect 32674 41964 32680 41976
rect 32732 41964 32738 42016
rect 34146 42004 34152 42016
rect 34107 41976 34152 42004
rect 34146 41964 34152 41976
rect 34204 41964 34210 42016
rect 37642 42004 37648 42016
rect 37603 41976 37648 42004
rect 37642 41964 37648 41976
rect 37700 41964 37706 42016
rect 38102 41964 38108 42016
rect 38160 42004 38166 42016
rect 38197 42007 38255 42013
rect 38197 42004 38209 42007
rect 38160 41976 38209 42004
rect 38160 41964 38166 41976
rect 38197 41973 38209 41976
rect 38243 42004 38255 42007
rect 38286 42004 38292 42016
rect 38243 41976 38292 42004
rect 38243 41973 38255 41976
rect 38197 41967 38255 41973
rect 38286 41964 38292 41976
rect 38344 41964 38350 42016
rect 42061 42007 42119 42013
rect 42061 41973 42073 42007
rect 42107 42004 42119 42007
rect 42334 42004 42340 42016
rect 42107 41976 42340 42004
rect 42107 41973 42119 41976
rect 42061 41967 42119 41973
rect 42334 41964 42340 41976
rect 42392 41964 42398 42016
rect 42444 42004 42472 42044
rect 44008 42004 44036 42180
rect 45189 42177 45201 42180
rect 45235 42208 45247 42211
rect 45278 42208 45284 42220
rect 45235 42180 45284 42208
rect 45235 42177 45247 42180
rect 45189 42171 45247 42177
rect 45278 42168 45284 42180
rect 45336 42168 45342 42220
rect 46934 42208 46940 42220
rect 46895 42180 46940 42208
rect 46934 42168 46940 42180
rect 46992 42168 46998 42220
rect 47213 42211 47271 42217
rect 47213 42177 47225 42211
rect 47259 42208 47271 42211
rect 47302 42208 47308 42220
rect 47259 42180 47308 42208
rect 47259 42177 47271 42180
rect 47213 42171 47271 42177
rect 47302 42168 47308 42180
rect 47360 42168 47366 42220
rect 47959 42217 47987 42316
rect 48958 42304 48964 42316
rect 49016 42304 49022 42356
rect 49050 42304 49056 42356
rect 49108 42344 49114 42356
rect 50249 42347 50307 42353
rect 50249 42344 50261 42347
rect 49108 42316 50261 42344
rect 49108 42304 49114 42316
rect 50249 42313 50261 42316
rect 50295 42344 50307 42347
rect 52454 42344 52460 42356
rect 50295 42316 52460 42344
rect 50295 42313 50307 42316
rect 50249 42307 50307 42313
rect 52454 42304 52460 42316
rect 52512 42304 52518 42356
rect 52638 42304 52644 42356
rect 52696 42344 52702 42356
rect 52696 42316 52960 42344
rect 52696 42304 52702 42316
rect 48130 42276 48136 42288
rect 48091 42248 48136 42276
rect 48130 42236 48136 42248
rect 48188 42236 48194 42288
rect 48682 42236 48688 42288
rect 48740 42276 48746 42288
rect 48866 42276 48872 42288
rect 48740 42248 48872 42276
rect 48740 42236 48746 42248
rect 48866 42236 48872 42248
rect 48924 42276 48930 42288
rect 48924 42248 52868 42276
rect 48924 42236 48930 42248
rect 47944 42211 48002 42217
rect 47944 42177 47956 42211
rect 47990 42177 48002 42211
rect 47944 42171 48002 42177
rect 48038 42168 48044 42220
rect 48096 42208 48102 42220
rect 48096 42180 48141 42208
rect 48096 42168 48102 42180
rect 48222 42168 48228 42220
rect 48280 42217 48286 42220
rect 49068 42217 49096 42248
rect 48280 42211 48319 42217
rect 48307 42177 48319 42211
rect 48280 42171 48319 42177
rect 48409 42211 48467 42217
rect 48409 42177 48421 42211
rect 48455 42177 48467 42211
rect 48409 42171 48467 42177
rect 49053 42211 49111 42217
rect 49053 42177 49065 42211
rect 49099 42177 49111 42211
rect 49234 42208 49240 42220
rect 49195 42180 49240 42208
rect 49053 42171 49111 42177
rect 48280 42168 48286 42171
rect 45094 42140 45100 42152
rect 45055 42112 45100 42140
rect 45094 42100 45100 42112
rect 45152 42100 45158 42152
rect 48424 42140 48452 42171
rect 49234 42168 49240 42180
rect 49292 42168 49298 42220
rect 49329 42211 49387 42217
rect 49329 42177 49341 42211
rect 49375 42177 49387 42211
rect 49329 42171 49387 42177
rect 49421 42211 49479 42217
rect 49421 42177 49433 42211
rect 49467 42208 49479 42211
rect 49602 42208 49608 42220
rect 49467 42180 49608 42208
rect 49467 42177 49479 42180
rect 49421 42171 49479 42177
rect 49344 42140 49372 42171
rect 49602 42168 49608 42180
rect 49660 42168 49666 42220
rect 49970 42168 49976 42220
rect 50028 42208 50034 42220
rect 50893 42211 50951 42217
rect 50893 42208 50905 42211
rect 50028 42180 50905 42208
rect 50028 42168 50034 42180
rect 50893 42177 50905 42180
rect 50939 42177 50951 42211
rect 50893 42171 50951 42177
rect 46952 42112 48452 42140
rect 48884 42112 49372 42140
rect 50985 42143 51043 42149
rect 46952 42081 46980 42112
rect 46937 42075 46995 42081
rect 46937 42041 46949 42075
rect 46983 42041 46995 42075
rect 48038 42072 48044 42084
rect 46937 42035 46995 42041
rect 47412 42044 48044 42072
rect 42444 41976 44036 42004
rect 44266 41964 44272 42016
rect 44324 42004 44330 42016
rect 44453 42007 44511 42013
rect 44453 42004 44465 42007
rect 44324 41976 44465 42004
rect 44324 41964 44330 41976
rect 44453 41973 44465 41976
rect 44499 42004 44511 42007
rect 47412 42004 47440 42044
rect 48038 42032 48044 42044
rect 48096 42072 48102 42084
rect 48096 42044 48314 42072
rect 48096 42032 48102 42044
rect 44499 41976 47440 42004
rect 44499 41973 44511 41976
rect 44453 41967 44511 41973
rect 47486 41964 47492 42016
rect 47544 42004 47550 42016
rect 47765 42007 47823 42013
rect 47765 42004 47777 42007
rect 47544 41976 47777 42004
rect 47544 41964 47550 41976
rect 47765 41973 47777 41976
rect 47811 41973 47823 42007
rect 48286 42004 48314 42044
rect 48406 42032 48412 42084
rect 48464 42072 48470 42084
rect 48884 42072 48912 42112
rect 50985 42109 50997 42143
rect 51031 42140 51043 42143
rect 51074 42140 51080 42152
rect 51031 42112 51080 42140
rect 51031 42109 51043 42112
rect 50985 42103 51043 42109
rect 51074 42100 51080 42112
rect 51132 42100 51138 42152
rect 51258 42140 51264 42152
rect 51219 42112 51264 42140
rect 51258 42100 51264 42112
rect 51316 42100 51322 42152
rect 52086 42100 52092 42152
rect 52144 42140 52150 42152
rect 52273 42143 52331 42149
rect 52273 42140 52285 42143
rect 52144 42112 52285 42140
rect 52144 42100 52150 42112
rect 52273 42109 52285 42112
rect 52319 42109 52331 42143
rect 52840 42140 52868 42248
rect 52932 42217 52960 42316
rect 53098 42304 53104 42356
rect 53156 42344 53162 42356
rect 53193 42347 53251 42353
rect 53193 42344 53205 42347
rect 53156 42316 53205 42344
rect 53156 42304 53162 42316
rect 53193 42313 53205 42316
rect 53239 42313 53251 42347
rect 54754 42344 54760 42356
rect 54715 42316 54760 42344
rect 53193 42307 53251 42313
rect 54754 42304 54760 42316
rect 54812 42304 54818 42356
rect 55122 42304 55128 42356
rect 55180 42344 55186 42356
rect 55769 42347 55827 42353
rect 55769 42344 55781 42347
rect 55180 42316 55781 42344
rect 55180 42304 55186 42316
rect 55769 42313 55781 42316
rect 55815 42344 55827 42347
rect 57330 42344 57336 42356
rect 55815 42316 57336 42344
rect 55815 42313 55827 42316
rect 55769 42307 55827 42313
rect 57330 42304 57336 42316
rect 57388 42304 57394 42356
rect 53650 42236 53656 42288
rect 53708 42276 53714 42288
rect 53708 42248 54616 42276
rect 53708 42236 53714 42248
rect 54588 42220 54616 42248
rect 55030 42236 55036 42288
rect 55088 42276 55094 42288
rect 55217 42279 55275 42285
rect 55217 42276 55229 42279
rect 55088 42248 55229 42276
rect 55088 42236 55094 42248
rect 55217 42245 55229 42248
rect 55263 42276 55275 42279
rect 56321 42279 56379 42285
rect 56321 42276 56333 42279
rect 55263 42248 56333 42276
rect 55263 42245 55275 42248
rect 55217 42239 55275 42245
rect 56321 42245 56333 42248
rect 56367 42245 56379 42279
rect 56321 42239 56379 42245
rect 52917 42211 52975 42217
rect 52917 42177 52929 42211
rect 52963 42177 52975 42211
rect 52917 42171 52975 42177
rect 53006 42168 53012 42220
rect 53064 42208 53070 42220
rect 53742 42208 53748 42220
rect 53064 42180 53748 42208
rect 53064 42168 53070 42180
rect 53742 42168 53748 42180
rect 53800 42168 53806 42220
rect 54110 42208 54116 42220
rect 54071 42180 54116 42208
rect 54110 42168 54116 42180
rect 54168 42168 54174 42220
rect 54294 42217 54300 42220
rect 54261 42211 54300 42217
rect 54261 42177 54273 42211
rect 54261 42171 54300 42177
rect 54294 42168 54300 42171
rect 54352 42168 54358 42220
rect 54389 42211 54447 42217
rect 54389 42177 54401 42211
rect 54435 42177 54447 42211
rect 54389 42171 54447 42177
rect 54481 42211 54539 42217
rect 54481 42177 54493 42211
rect 54527 42177 54539 42211
rect 54481 42171 54539 42177
rect 53190 42140 53196 42152
rect 52840 42112 53196 42140
rect 52273 42103 52331 42109
rect 53190 42100 53196 42112
rect 53248 42140 53254 42152
rect 53374 42140 53380 42152
rect 53248 42112 53380 42140
rect 53248 42100 53254 42112
rect 53374 42100 53380 42112
rect 53432 42100 53438 42152
rect 53926 42100 53932 42152
rect 53984 42140 53990 42152
rect 54404 42140 54432 42171
rect 53984 42112 54432 42140
rect 54496 42140 54524 42171
rect 54570 42168 54576 42220
rect 54628 42217 54634 42220
rect 54628 42208 54636 42217
rect 54628 42180 54673 42208
rect 54628 42171 54636 42180
rect 54628 42168 54634 42171
rect 55030 42140 55036 42152
rect 54496 42112 55036 42140
rect 53984 42100 53990 42112
rect 55030 42100 55036 42112
rect 55088 42100 55094 42152
rect 48464 42044 48912 42072
rect 48464 42032 48470 42044
rect 49418 42032 49424 42084
rect 49476 42072 49482 42084
rect 51718 42072 51724 42084
rect 49476 42044 51724 42072
rect 49476 42032 49482 42044
rect 51718 42032 51724 42044
rect 51776 42032 51782 42084
rect 52196 42044 52592 42072
rect 52196 42016 52224 42044
rect 49050 42004 49056 42016
rect 48286 41976 49056 42004
rect 47765 41967 47823 41973
rect 49050 41964 49056 41976
rect 49108 41964 49114 42016
rect 49694 42004 49700 42016
rect 49655 41976 49700 42004
rect 49694 41964 49700 41976
rect 49752 41964 49758 42016
rect 51813 42007 51871 42013
rect 51813 41973 51825 42007
rect 51859 42004 51871 42007
rect 52178 42004 52184 42016
rect 51859 41976 52184 42004
rect 51859 41973 51871 41976
rect 51813 41967 51871 41973
rect 52178 41964 52184 41976
rect 52236 41964 52242 42016
rect 52564 42004 52592 42044
rect 53098 42004 53104 42016
rect 52564 41976 53104 42004
rect 53098 41964 53104 41976
rect 53156 41964 53162 42016
rect 54018 41964 54024 42016
rect 54076 42004 54082 42016
rect 54386 42004 54392 42016
rect 54076 41976 54392 42004
rect 54076 41964 54082 41976
rect 54386 41964 54392 41976
rect 54444 41964 54450 42016
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 33686 41800 33692 41812
rect 33647 41772 33692 41800
rect 33686 41760 33692 41772
rect 33744 41760 33750 41812
rect 36633 41803 36691 41809
rect 36633 41769 36645 41803
rect 36679 41800 36691 41803
rect 36722 41800 36728 41812
rect 36679 41772 36728 41800
rect 36679 41769 36691 41772
rect 36633 41763 36691 41769
rect 36722 41760 36728 41772
rect 36780 41760 36786 41812
rect 40770 41800 40776 41812
rect 40731 41772 40776 41800
rect 40770 41760 40776 41772
rect 40828 41760 40834 41812
rect 45094 41800 45100 41812
rect 41386 41772 45100 41800
rect 31018 41732 31024 41744
rect 30979 41704 31024 41732
rect 31018 41692 31024 41704
rect 31076 41692 31082 41744
rect 41386 41732 41414 41772
rect 45094 41760 45100 41772
rect 45152 41800 45158 41812
rect 45152 41772 45508 41800
rect 45152 41760 45158 41772
rect 36004 41704 41414 41732
rect 28902 41664 28908 41676
rect 28863 41636 28908 41664
rect 28902 41624 28908 41636
rect 28960 41624 28966 41676
rect 29181 41667 29239 41673
rect 29181 41633 29193 41667
rect 29227 41664 29239 41667
rect 30009 41667 30067 41673
rect 30009 41664 30021 41667
rect 29227 41636 30021 41664
rect 29227 41633 29239 41636
rect 29181 41627 29239 41633
rect 30009 41633 30021 41636
rect 30055 41633 30067 41667
rect 30009 41627 30067 41633
rect 30650 41624 30656 41676
rect 30708 41664 30714 41676
rect 31846 41664 31852 41676
rect 30708 41636 30972 41664
rect 31807 41636 31852 41664
rect 30708 41624 30714 41636
rect 28813 41599 28871 41605
rect 28813 41565 28825 41599
rect 28859 41596 28871 41599
rect 29270 41596 29276 41608
rect 28859 41568 29276 41596
rect 28859 41565 28871 41568
rect 28813 41559 28871 41565
rect 29270 41556 29276 41568
rect 29328 41556 29334 41608
rect 30101 41599 30159 41605
rect 30101 41565 30113 41599
rect 30147 41596 30159 41599
rect 30834 41596 30840 41608
rect 30147 41568 30840 41596
rect 30147 41565 30159 41568
rect 30101 41559 30159 41565
rect 30834 41556 30840 41568
rect 30892 41556 30898 41608
rect 30944 41605 30972 41636
rect 31846 41624 31852 41636
rect 31904 41624 31910 41676
rect 33318 41664 33324 41676
rect 33279 41636 33324 41664
rect 33318 41624 33324 41636
rect 33376 41624 33382 41676
rect 34698 41624 34704 41676
rect 34756 41664 34762 41676
rect 36004 41673 36032 41704
rect 42886 41692 42892 41744
rect 42944 41692 42950 41744
rect 42981 41735 43039 41741
rect 42981 41701 42993 41735
rect 43027 41701 43039 41735
rect 42981 41695 43039 41701
rect 35989 41667 36047 41673
rect 34756 41636 35296 41664
rect 34756 41624 34762 41636
rect 30929 41599 30987 41605
rect 30929 41565 30941 41599
rect 30975 41565 30987 41599
rect 30929 41559 30987 41565
rect 31757 41599 31815 41605
rect 31757 41565 31769 41599
rect 31803 41596 31815 41599
rect 31938 41596 31944 41608
rect 31803 41568 31944 41596
rect 31803 41565 31815 41568
rect 31757 41559 31815 41565
rect 31938 41556 31944 41568
rect 31996 41556 32002 41608
rect 32214 41596 32220 41608
rect 32175 41568 32220 41596
rect 32214 41556 32220 41568
rect 32272 41556 32278 41608
rect 32766 41596 32772 41608
rect 32727 41568 32772 41596
rect 32766 41556 32772 41568
rect 32824 41556 32830 41608
rect 33413 41599 33471 41605
rect 33413 41565 33425 41599
rect 33459 41565 33471 41599
rect 34974 41596 34980 41608
rect 34935 41568 34980 41596
rect 33413 41559 33471 41565
rect 32858 41528 32864 41540
rect 30484 41500 32864 41528
rect 30484 41469 30512 41500
rect 32858 41488 32864 41500
rect 32916 41528 32922 41540
rect 33428 41528 33456 41559
rect 34974 41556 34980 41568
rect 35032 41556 35038 41608
rect 35161 41599 35219 41605
rect 35161 41565 35173 41599
rect 35207 41565 35219 41599
rect 35268 41596 35296 41636
rect 35989 41633 36001 41667
rect 36035 41633 36047 41667
rect 35989 41627 36047 41633
rect 37550 41624 37556 41676
rect 37608 41664 37614 41676
rect 38010 41664 38016 41676
rect 37608 41636 38016 41664
rect 37608 41624 37614 41636
rect 38010 41624 38016 41636
rect 38068 41624 38074 41676
rect 38654 41664 38660 41676
rect 38615 41636 38660 41664
rect 38654 41624 38660 41636
rect 38712 41624 38718 41676
rect 40770 41664 40776 41676
rect 40509 41636 40776 41664
rect 36449 41599 36507 41605
rect 36449 41596 36461 41599
rect 35268 41568 36461 41596
rect 35161 41559 35219 41565
rect 36449 41565 36461 41568
rect 36495 41565 36507 41599
rect 36449 41559 36507 41565
rect 37461 41599 37519 41605
rect 37461 41565 37473 41599
rect 37507 41596 37519 41599
rect 37734 41596 37740 41608
rect 37507 41568 37740 41596
rect 37507 41565 37519 41568
rect 37461 41559 37519 41565
rect 32916 41500 33456 41528
rect 32916 41488 32922 41500
rect 33962 41488 33968 41540
rect 34020 41528 34026 41540
rect 35176 41528 35204 41559
rect 37734 41556 37740 41568
rect 37792 41556 37798 41608
rect 37829 41599 37887 41605
rect 37829 41565 37841 41599
rect 37875 41596 37887 41599
rect 37918 41596 37924 41608
rect 37875 41568 37924 41596
rect 37875 41565 37887 41568
rect 37829 41559 37887 41565
rect 37918 41556 37924 41568
rect 37976 41556 37982 41608
rect 38102 41596 38108 41608
rect 38063 41568 38108 41596
rect 38102 41556 38108 41568
rect 38160 41556 38166 41608
rect 38749 41599 38807 41605
rect 38749 41565 38761 41599
rect 38795 41596 38807 41599
rect 39206 41596 39212 41608
rect 38795 41568 39212 41596
rect 38795 41565 38807 41568
rect 38749 41559 38807 41565
rect 39206 41556 39212 41568
rect 39264 41556 39270 41608
rect 40126 41596 40132 41608
rect 40087 41568 40132 41596
rect 40126 41556 40132 41568
rect 40184 41556 40190 41608
rect 40218 41556 40224 41608
rect 40276 41605 40282 41608
rect 40509 41605 40537 41636
rect 40770 41624 40776 41636
rect 40828 41664 40834 41676
rect 41874 41664 41880 41676
rect 40828 41636 41880 41664
rect 40828 41624 40834 41636
rect 41874 41624 41880 41636
rect 41932 41664 41938 41676
rect 42904 41664 42932 41692
rect 41932 41636 42473 41664
rect 41932 41624 41938 41636
rect 40678 41605 40684 41608
rect 40276 41599 40307 41605
rect 40295 41596 40307 41599
rect 40494 41599 40552 41605
rect 40295 41568 40369 41596
rect 40295 41565 40307 41568
rect 40276 41559 40307 41565
rect 40494 41565 40506 41599
rect 40540 41565 40552 41599
rect 40494 41559 40552 41565
rect 40633 41599 40684 41605
rect 40633 41565 40645 41599
rect 40679 41565 40684 41599
rect 40633 41559 40684 41565
rect 40276 41556 40282 41559
rect 40678 41556 40684 41559
rect 40736 41596 40742 41608
rect 40954 41596 40960 41608
rect 40736 41568 40960 41596
rect 40736 41556 40742 41568
rect 40954 41556 40960 41568
rect 41012 41556 41018 41608
rect 41322 41596 41328 41608
rect 41283 41568 41328 41596
rect 41322 41556 41328 41568
rect 41380 41556 41386 41608
rect 42334 41596 42340 41608
rect 42295 41568 42340 41596
rect 42334 41556 42340 41568
rect 42392 41556 42398 41608
rect 42445 41605 42473 41636
rect 42628 41636 42932 41664
rect 42430 41599 42488 41605
rect 42430 41565 42442 41599
rect 42476 41596 42488 41599
rect 42518 41596 42524 41608
rect 42476 41568 42524 41596
rect 42476 41565 42488 41568
rect 42430 41559 42488 41565
rect 42518 41556 42524 41568
rect 42576 41556 42582 41608
rect 42628 41605 42656 41636
rect 42613 41599 42671 41605
rect 42613 41565 42625 41599
rect 42659 41565 42671 41599
rect 42613 41559 42671 41565
rect 42802 41599 42860 41605
rect 42802 41565 42814 41599
rect 42848 41596 42860 41599
rect 42996 41596 43024 41695
rect 43898 41664 43904 41676
rect 43859 41636 43904 41664
rect 43898 41624 43904 41636
rect 43956 41624 43962 41676
rect 44177 41667 44235 41673
rect 44177 41633 44189 41667
rect 44223 41664 44235 41667
rect 45373 41667 45431 41673
rect 45373 41664 45385 41667
rect 44223 41636 45385 41664
rect 44223 41633 44235 41636
rect 44177 41627 44235 41633
rect 45373 41633 45385 41636
rect 45419 41633 45431 41667
rect 45373 41627 45431 41633
rect 45480 41605 45508 41772
rect 47578 41760 47584 41812
rect 47636 41800 47642 41812
rect 48130 41800 48136 41812
rect 47636 41772 48136 41800
rect 47636 41760 47642 41772
rect 48130 41760 48136 41772
rect 48188 41760 48194 41812
rect 48593 41803 48651 41809
rect 48593 41769 48605 41803
rect 48639 41800 48651 41803
rect 49050 41800 49056 41812
rect 48639 41772 49056 41800
rect 48639 41769 48651 41772
rect 48593 41763 48651 41769
rect 49050 41760 49056 41772
rect 49108 41760 49114 41812
rect 49145 41803 49203 41809
rect 49145 41769 49157 41803
rect 49191 41800 49203 41803
rect 49234 41800 49240 41812
rect 49191 41772 49240 41800
rect 49191 41769 49203 41772
rect 49145 41763 49203 41769
rect 49234 41760 49240 41772
rect 49292 41760 49298 41812
rect 51074 41800 51080 41812
rect 49533 41772 51080 41800
rect 49533 41732 49561 41772
rect 51074 41760 51080 41772
rect 51132 41760 51138 41812
rect 54665 41803 54723 41809
rect 54665 41800 54677 41803
rect 52472 41772 54677 41800
rect 51902 41732 51908 41744
rect 46308 41704 49561 41732
rect 49625 41704 51908 41732
rect 46308 41673 46336 41704
rect 46293 41667 46351 41673
rect 46293 41633 46305 41667
rect 46339 41633 46351 41667
rect 47486 41664 47492 41676
rect 47447 41636 47492 41664
rect 46293 41627 46351 41633
rect 47486 41624 47492 41636
rect 47544 41624 47550 41676
rect 43809 41599 43867 41605
rect 43809 41596 43821 41599
rect 42848 41568 42932 41596
rect 42996 41568 43821 41596
rect 42848 41565 42860 41568
rect 42802 41559 42860 41565
rect 34020 41500 35204 41528
rect 34020 41488 34026 41500
rect 37182 41488 37188 41540
rect 37240 41528 37246 41540
rect 40236 41528 40264 41556
rect 40402 41528 40408 41540
rect 37240 41500 40264 41528
rect 40363 41500 40408 41528
rect 37240 41488 37246 41500
rect 40402 41488 40408 41500
rect 40460 41488 40466 41540
rect 30469 41463 30527 41469
rect 30469 41429 30481 41463
rect 30515 41429 30527 41463
rect 30469 41423 30527 41429
rect 37642 41420 37648 41472
rect 37700 41460 37706 41472
rect 40696 41460 40724 41556
rect 37700 41432 40724 41460
rect 41340 41460 41368 41556
rect 41693 41531 41751 41537
rect 41693 41497 41705 41531
rect 41739 41528 41751 41531
rect 42242 41528 42248 41540
rect 41739 41500 42248 41528
rect 41739 41497 41751 41500
rect 41693 41491 41751 41497
rect 42242 41488 42248 41500
rect 42300 41488 42306 41540
rect 42705 41531 42763 41537
rect 42705 41497 42717 41531
rect 42751 41497 42763 41531
rect 42904 41528 42932 41568
rect 43809 41565 43821 41568
rect 43855 41565 43867 41599
rect 43809 41559 43867 41565
rect 45465 41599 45523 41605
rect 45465 41565 45477 41599
rect 45511 41565 45523 41599
rect 47394 41596 47400 41608
rect 47355 41568 47400 41596
rect 45465 41559 45523 41565
rect 47394 41556 47400 41568
rect 47452 41556 47458 41608
rect 48314 41596 48320 41608
rect 48275 41568 48320 41596
rect 48314 41556 48320 41568
rect 48372 41556 48378 41608
rect 49050 41556 49056 41608
rect 49108 41596 49114 41608
rect 49518 41599 49576 41605
rect 49518 41596 49530 41599
rect 49108 41568 49530 41596
rect 49108 41556 49114 41568
rect 49518 41565 49530 41568
rect 49564 41596 49576 41599
rect 49625 41596 49653 41704
rect 51902 41692 51908 41704
rect 51960 41692 51966 41744
rect 52086 41692 52092 41744
rect 52144 41732 52150 41744
rect 52472 41732 52500 41772
rect 54665 41769 54677 41772
rect 54711 41769 54723 41803
rect 54665 41763 54723 41769
rect 52144 41704 52500 41732
rect 52144 41692 52150 41704
rect 49694 41624 49700 41676
rect 49752 41664 49758 41676
rect 50433 41667 50491 41673
rect 50433 41664 50445 41667
rect 49752 41636 50445 41664
rect 49752 41624 49758 41636
rect 50433 41633 50445 41636
rect 50479 41633 50491 41667
rect 50433 41627 50491 41633
rect 51534 41624 51540 41676
rect 51592 41664 51598 41676
rect 51592 41636 52224 41664
rect 51592 41624 51598 41636
rect 52196 41608 52224 41636
rect 50522 41596 50528 41608
rect 49564 41568 49653 41596
rect 50483 41568 50528 41596
rect 49564 41565 49576 41568
rect 49518 41559 49576 41565
rect 50522 41556 50528 41568
rect 50580 41556 50586 41608
rect 51166 41556 51172 41608
rect 51224 41596 51230 41608
rect 52089 41599 52147 41605
rect 52089 41596 52101 41599
rect 51224 41568 52101 41596
rect 51224 41556 51230 41568
rect 52089 41565 52101 41568
rect 52135 41565 52147 41599
rect 52089 41559 52147 41565
rect 52178 41556 52184 41608
rect 52236 41596 52242 41608
rect 52472 41605 52500 41704
rect 52733 41735 52791 41741
rect 52733 41701 52745 41735
rect 52779 41732 52791 41735
rect 52779 41704 56180 41732
rect 52779 41701 52791 41704
rect 52733 41695 52791 41701
rect 52638 41624 52644 41676
rect 52696 41664 52702 41676
rect 52696 41636 52960 41664
rect 52696 41624 52702 41636
rect 52457 41599 52515 41605
rect 52236 41568 52281 41596
rect 52236 41556 52242 41568
rect 52457 41565 52469 41599
rect 52503 41565 52515 41599
rect 52457 41559 52515 41565
rect 52554 41599 52612 41605
rect 52554 41565 52566 41599
rect 52600 41596 52612 41599
rect 52822 41596 52828 41608
rect 52600 41568 52828 41596
rect 52600 41565 52612 41568
rect 52554 41559 52612 41565
rect 52822 41556 52828 41568
rect 52880 41556 52886 41608
rect 52932 41596 52960 41636
rect 53098 41624 53104 41676
rect 53156 41664 53162 41676
rect 53193 41667 53251 41673
rect 53193 41664 53205 41667
rect 53156 41636 53205 41664
rect 53156 41624 53162 41636
rect 53193 41633 53205 41636
rect 53239 41664 53251 41667
rect 53558 41664 53564 41676
rect 53239 41636 53564 41664
rect 53239 41633 53251 41636
rect 53193 41627 53251 41633
rect 53558 41624 53564 41636
rect 53616 41624 53622 41676
rect 54018 41664 54024 41676
rect 53979 41636 54024 41664
rect 54018 41624 54024 41636
rect 54076 41624 54082 41676
rect 56152 41673 56180 41704
rect 56137 41667 56195 41673
rect 56137 41633 56149 41667
rect 56183 41633 56195 41667
rect 56137 41627 56195 41633
rect 57057 41667 57115 41673
rect 57057 41633 57069 41667
rect 57103 41664 57115 41667
rect 57238 41664 57244 41676
rect 57103 41636 57244 41664
rect 57103 41633 57115 41636
rect 57057 41627 57115 41633
rect 57238 41624 57244 41636
rect 57296 41664 57302 41676
rect 57422 41664 57428 41676
rect 57296 41636 57428 41664
rect 57296 41624 57302 41636
rect 57422 41624 57428 41636
rect 57480 41624 57486 41676
rect 53745 41599 53803 41605
rect 53745 41596 53757 41599
rect 52932 41568 53757 41596
rect 53745 41565 53757 41568
rect 53791 41565 53803 41599
rect 53926 41596 53932 41608
rect 53887 41568 53932 41596
rect 53745 41559 53803 41565
rect 53926 41556 53932 41568
rect 53984 41556 53990 41608
rect 54118 41599 54176 41605
rect 54118 41565 54130 41599
rect 54164 41565 54176 41599
rect 56226 41596 56232 41608
rect 56187 41568 56232 41596
rect 54118 41559 54176 41565
rect 43070 41528 43076 41540
rect 42904 41500 43076 41528
rect 42705 41491 42763 41497
rect 42720 41460 42748 41491
rect 43070 41488 43076 41500
rect 43128 41488 43134 41540
rect 48774 41488 48780 41540
rect 48832 41528 48838 41540
rect 49145 41531 49203 41537
rect 49145 41528 49157 41531
rect 48832 41500 49157 41528
rect 48832 41488 48838 41500
rect 49145 41497 49157 41500
rect 49191 41528 49203 41531
rect 49234 41528 49240 41540
rect 49191 41500 49240 41528
rect 49191 41497 49203 41500
rect 49145 41491 49203 41497
rect 49234 41488 49240 41500
rect 49292 41488 49298 41540
rect 49329 41531 49387 41537
rect 49329 41497 49341 41531
rect 49375 41497 49387 41531
rect 49329 41491 49387 41497
rect 49421 41531 49479 41537
rect 49421 41497 49433 41531
rect 49467 41528 49479 41531
rect 49602 41528 49608 41540
rect 49467 41500 49608 41528
rect 49467 41497 49479 41500
rect 49421 41491 49479 41497
rect 43714 41460 43720 41472
rect 41340 41432 43720 41460
rect 37700 41420 37706 41432
rect 43714 41420 43720 41432
rect 43772 41420 43778 41472
rect 47765 41463 47823 41469
rect 47765 41429 47777 41463
rect 47811 41460 47823 41463
rect 47946 41460 47952 41472
rect 47811 41432 47952 41460
rect 47811 41429 47823 41432
rect 47765 41423 47823 41429
rect 47946 41420 47952 41432
rect 48004 41420 48010 41472
rect 49344 41460 49372 41491
rect 49602 41488 49608 41500
rect 49660 41488 49666 41540
rect 49712 41500 52224 41528
rect 49712 41460 49740 41500
rect 49344 41432 49740 41460
rect 49786 41420 49792 41472
rect 49844 41460 49850 41472
rect 49970 41460 49976 41472
rect 49844 41432 49976 41460
rect 49844 41420 49850 41432
rect 49970 41420 49976 41432
rect 50028 41420 50034 41472
rect 50890 41460 50896 41472
rect 50851 41432 50896 41460
rect 50890 41420 50896 41432
rect 50948 41420 50954 41472
rect 50982 41420 50988 41472
rect 51040 41460 51046 41472
rect 51353 41463 51411 41469
rect 51353 41460 51365 41463
rect 51040 41432 51365 41460
rect 51040 41420 51046 41432
rect 51353 41429 51365 41432
rect 51399 41460 51411 41463
rect 51718 41460 51724 41472
rect 51399 41432 51724 41460
rect 51399 41429 51411 41432
rect 51353 41423 51411 41429
rect 51718 41420 51724 41432
rect 51776 41460 51782 41472
rect 51994 41460 52000 41472
rect 51776 41432 52000 41460
rect 51776 41420 51782 41432
rect 51994 41420 52000 41432
rect 52052 41420 52058 41472
rect 52196 41460 52224 41500
rect 52270 41488 52276 41540
rect 52328 41528 52334 41540
rect 52365 41531 52423 41537
rect 52365 41528 52377 41531
rect 52328 41500 52377 41528
rect 52328 41488 52334 41500
rect 52365 41497 52377 41500
rect 52411 41497 52423 41531
rect 54021 41531 54079 41537
rect 52365 41491 52423 41497
rect 52564 41500 53604 41528
rect 52564 41460 52592 41500
rect 52196 41432 52592 41460
rect 53576 41460 53604 41500
rect 54021 41497 54033 41531
rect 54067 41497 54079 41531
rect 54133 41528 54161 41559
rect 56226 41556 56232 41568
rect 56284 41556 56290 41608
rect 54386 41528 54392 41540
rect 54133 41500 54392 41528
rect 54021 41491 54079 41497
rect 53834 41460 53840 41472
rect 53576 41432 53840 41460
rect 53834 41420 53840 41432
rect 53892 41420 53898 41472
rect 54036 41460 54064 41491
rect 54386 41488 54392 41500
rect 54444 41488 54450 41540
rect 54294 41460 54300 41472
rect 54036 41432 54300 41460
rect 54294 41420 54300 41432
rect 54352 41420 54358 41472
rect 54478 41420 54484 41472
rect 54536 41460 54542 41472
rect 55030 41460 55036 41472
rect 54536 41432 55036 41460
rect 54536 41420 54542 41432
rect 55030 41420 55036 41432
rect 55088 41420 55094 41472
rect 1104 41370 58880 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 35594 41370
rect 35646 41318 35658 41370
rect 35710 41318 35722 41370
rect 35774 41318 35786 41370
rect 35838 41318 35850 41370
rect 35902 41318 58880 41370
rect 1104 41296 58880 41318
rect 32861 41259 32919 41265
rect 32861 41225 32873 41259
rect 32907 41225 32919 41259
rect 32861 41219 32919 41225
rect 33873 41259 33931 41265
rect 33873 41225 33885 41259
rect 33919 41256 33931 41259
rect 34974 41256 34980 41268
rect 33919 41228 34980 41256
rect 33919 41225 33931 41228
rect 33873 41219 33931 41225
rect 32306 41080 32312 41132
rect 32364 41120 32370 41132
rect 32493 41123 32551 41129
rect 32493 41120 32505 41123
rect 32364 41092 32505 41120
rect 32364 41080 32370 41092
rect 32493 41089 32505 41092
rect 32539 41089 32551 41123
rect 32876 41120 32904 41219
rect 34974 41216 34980 41228
rect 35032 41216 35038 41268
rect 36541 41259 36599 41265
rect 36541 41225 36553 41259
rect 36587 41256 36599 41259
rect 36630 41256 36636 41268
rect 36587 41228 36636 41256
rect 36587 41225 36599 41228
rect 36541 41219 36599 41225
rect 36630 41216 36636 41228
rect 36688 41216 36694 41268
rect 37458 41216 37464 41268
rect 37516 41256 37522 41268
rect 37516 41228 37872 41256
rect 37516 41216 37522 41228
rect 34790 41148 34796 41200
rect 34848 41188 34854 41200
rect 35621 41191 35679 41197
rect 35621 41188 35633 41191
rect 34848 41160 35633 41188
rect 34848 41148 34854 41160
rect 35621 41157 35633 41160
rect 35667 41188 35679 41191
rect 37844 41188 37872 41228
rect 38378 41216 38384 41268
rect 38436 41256 38442 41268
rect 38436 41228 38516 41256
rect 38436 41216 38442 41228
rect 38102 41188 38108 41200
rect 35667 41160 36400 41188
rect 35667 41157 35679 41160
rect 35621 41151 35679 41157
rect 33318 41120 33324 41132
rect 32876 41092 33324 41120
rect 32493 41083 32551 41089
rect 33318 41080 33324 41092
rect 33376 41120 33382 41132
rect 35434 41129 35440 41132
rect 33505 41123 33563 41129
rect 33505 41120 33517 41123
rect 33376 41092 33517 41120
rect 33376 41080 33382 41092
rect 33505 41089 33517 41092
rect 33551 41089 33563 41123
rect 35432 41120 35440 41129
rect 35395 41092 35440 41120
rect 33505 41083 33563 41089
rect 35432 41083 35440 41092
rect 35434 41080 35440 41083
rect 35492 41080 35498 41132
rect 35526 41080 35532 41132
rect 35584 41120 35590 41132
rect 35802 41120 35808 41132
rect 35584 41092 35629 41120
rect 35763 41092 35808 41120
rect 35584 41080 35590 41092
rect 35802 41080 35808 41092
rect 35860 41080 35866 41132
rect 35894 41080 35900 41132
rect 35952 41120 35958 41132
rect 36372 41129 36400 41160
rect 37844 41160 38108 41188
rect 36357 41123 36415 41129
rect 35952 41092 35997 41120
rect 35952 41080 35958 41092
rect 36357 41089 36369 41123
rect 36403 41089 36415 41123
rect 36357 41083 36415 41089
rect 37274 41080 37280 41132
rect 37332 41120 37338 41132
rect 37461 41123 37519 41129
rect 37461 41120 37473 41123
rect 37332 41092 37473 41120
rect 37332 41080 37338 41092
rect 37461 41089 37473 41092
rect 37507 41089 37519 41123
rect 37461 41083 37519 41089
rect 37550 41080 37556 41132
rect 37608 41120 37614 41132
rect 37737 41123 37795 41129
rect 37608 41092 37653 41120
rect 37608 41080 37614 41092
rect 37737 41089 37749 41123
rect 37783 41120 37795 41123
rect 37844 41120 37872 41160
rect 38102 41148 38108 41160
rect 38160 41148 38166 41200
rect 38488 41197 38516 41228
rect 38562 41216 38568 41268
rect 38620 41216 38626 41268
rect 38841 41259 38899 41265
rect 38841 41225 38853 41259
rect 38887 41256 38899 41259
rect 38930 41256 38936 41268
rect 38887 41228 38936 41256
rect 38887 41225 38899 41228
rect 38841 41219 38899 41225
rect 38930 41216 38936 41228
rect 38988 41216 38994 41268
rect 40681 41259 40739 41265
rect 40681 41256 40693 41259
rect 39776 41228 40693 41256
rect 38473 41191 38531 41197
rect 38473 41157 38485 41191
rect 38519 41157 38531 41191
rect 38580 41188 38608 41216
rect 39776 41188 39804 41228
rect 40681 41225 40693 41228
rect 40727 41256 40739 41259
rect 44266 41256 44272 41268
rect 40727 41228 44272 41256
rect 40727 41225 40739 41228
rect 40681 41219 40739 41225
rect 44266 41216 44272 41228
rect 44324 41216 44330 41268
rect 47854 41256 47860 41268
rect 47815 41228 47860 41256
rect 47854 41216 47860 41228
rect 47912 41256 47918 41268
rect 48222 41256 48228 41268
rect 47912 41228 48228 41256
rect 47912 41216 47918 41228
rect 48222 41216 48228 41228
rect 48280 41216 48286 41268
rect 49234 41256 49240 41268
rect 49195 41228 49240 41256
rect 49234 41216 49240 41228
rect 49292 41216 49298 41268
rect 50246 41216 50252 41268
rect 50304 41256 50310 41268
rect 50893 41259 50951 41265
rect 50893 41256 50905 41259
rect 50304 41228 50905 41256
rect 50304 41216 50310 41228
rect 50893 41225 50905 41228
rect 50939 41225 50951 41259
rect 50893 41219 50951 41225
rect 51074 41216 51080 41268
rect 51132 41256 51138 41268
rect 55585 41259 55643 41265
rect 51132 41228 55260 41256
rect 51132 41216 51138 41228
rect 41877 41191 41935 41197
rect 41877 41188 41889 41191
rect 38580 41160 39804 41188
rect 41386 41160 41889 41188
rect 38473 41151 38531 41157
rect 37783 41092 37872 41120
rect 37783 41089 37795 41092
rect 37737 41083 37795 41089
rect 37918 41080 37924 41132
rect 37976 41120 37982 41132
rect 38378 41129 38384 41132
rect 38197 41123 38255 41129
rect 38197 41120 38209 41123
rect 37976 41092 38209 41120
rect 37976 41080 37982 41092
rect 38197 41089 38209 41092
rect 38243 41089 38255 41123
rect 38197 41083 38255 41089
rect 38335 41123 38384 41129
rect 38335 41089 38347 41123
rect 38381 41089 38384 41123
rect 38335 41083 38384 41089
rect 38378 41080 38384 41083
rect 38436 41080 38442 41132
rect 38608 41129 38614 41132
rect 38594 41123 38614 41129
rect 38594 41089 38606 41123
rect 38594 41083 38614 41089
rect 38608 41080 38614 41083
rect 38666 41080 38672 41132
rect 38746 41129 38752 41132
rect 38703 41123 38752 41129
rect 38703 41089 38715 41123
rect 38749 41089 38752 41123
rect 38703 41083 38752 41089
rect 38746 41080 38752 41083
rect 38804 41080 38810 41132
rect 39853 41123 39911 41129
rect 39853 41120 39865 41123
rect 39776 41092 39865 41120
rect 29086 41012 29092 41064
rect 29144 41052 29150 41064
rect 32401 41055 32459 41061
rect 32401 41052 32413 41055
rect 29144 41024 32413 41052
rect 29144 41012 29150 41024
rect 32401 41021 32413 41024
rect 32447 41021 32459 41055
rect 32401 41015 32459 41021
rect 33597 41055 33655 41061
rect 33597 41021 33609 41055
rect 33643 41021 33655 41055
rect 39776 41052 39804 41092
rect 39853 41089 39865 41092
rect 39899 41120 39911 41123
rect 40678 41120 40684 41132
rect 39899 41092 40684 41120
rect 39899 41089 39911 41092
rect 39853 41083 39911 41089
rect 40678 41080 40684 41092
rect 40736 41080 40742 41132
rect 33597 41015 33655 41021
rect 38626 41024 39804 41052
rect 40129 41055 40187 41061
rect 33612 40984 33640 41015
rect 38626 40996 38654 41024
rect 40129 41021 40141 41055
rect 40175 41021 40187 41055
rect 40129 41015 40187 41021
rect 35253 40987 35311 40993
rect 35253 40984 35265 40987
rect 33612 40956 35265 40984
rect 35253 40953 35265 40956
rect 35299 40953 35311 40987
rect 35253 40947 35311 40953
rect 35434 40944 35440 40996
rect 35492 40984 35498 40996
rect 35986 40984 35992 40996
rect 35492 40956 35992 40984
rect 35492 40944 35498 40956
rect 35986 40944 35992 40956
rect 36044 40944 36050 40996
rect 37734 40984 37740 40996
rect 37695 40956 37740 40984
rect 37734 40944 37740 40956
rect 37792 40944 37798 40996
rect 38562 40944 38568 40996
rect 38620 40956 38654 40996
rect 38620 40944 38626 40956
rect 39482 40944 39488 40996
rect 39540 40984 39546 40996
rect 40144 40984 40172 41015
rect 39540 40956 40172 40984
rect 39540 40944 39546 40956
rect 40770 40944 40776 40996
rect 40828 40984 40834 40996
rect 41386 40984 41414 41160
rect 41877 41157 41889 41160
rect 41923 41188 41935 41191
rect 42334 41188 42340 41200
rect 41923 41160 42340 41188
rect 41923 41157 41935 41160
rect 41877 41151 41935 41157
rect 42334 41148 42340 41160
rect 42392 41148 42398 41200
rect 42518 41148 42524 41200
rect 42576 41188 42582 41200
rect 42981 41191 43039 41197
rect 42981 41188 42993 41191
rect 42576 41160 42993 41188
rect 42576 41148 42582 41160
rect 42981 41157 42993 41160
rect 43027 41157 43039 41191
rect 43990 41188 43996 41200
rect 42981 41151 43039 41157
rect 43134 41160 43996 41188
rect 43134 41132 43162 41160
rect 43990 41148 43996 41160
rect 44048 41148 44054 41200
rect 47213 41191 47271 41197
rect 47213 41157 47225 41191
rect 47259 41188 47271 41191
rect 47259 41160 50752 41188
rect 47259 41157 47271 41160
rect 47213 41151 47271 41157
rect 41690 41080 41696 41132
rect 41748 41120 41754 41132
rect 41785 41123 41843 41129
rect 41785 41120 41797 41123
rect 41748 41092 41797 41120
rect 41748 41080 41754 41092
rect 41785 41089 41797 41092
rect 41831 41089 41843 41123
rect 41785 41083 41843 41089
rect 41966 41080 41972 41132
rect 42024 41120 42030 41132
rect 43134 41129 43168 41132
rect 42061 41123 42119 41129
rect 42061 41120 42073 41123
rect 42024 41092 42073 41120
rect 42024 41080 42030 41092
rect 42061 41089 42073 41092
rect 42107 41089 42119 41123
rect 42061 41083 42119 41089
rect 42613 41123 42671 41129
rect 42613 41089 42625 41123
rect 42659 41089 42671 41123
rect 42613 41083 42671 41089
rect 42706 41123 42764 41129
rect 42706 41089 42718 41123
rect 42752 41089 42764 41123
rect 42706 41083 42764 41089
rect 42889 41123 42947 41129
rect 42889 41089 42901 41123
rect 42935 41089 42947 41123
rect 42889 41083 42947 41089
rect 43119 41123 43168 41129
rect 43119 41089 43131 41123
rect 43165 41089 43168 41123
rect 43119 41083 43168 41089
rect 42628 41052 42656 41083
rect 42076 41024 42656 41052
rect 42076 40993 42104 41024
rect 40828 40956 41414 40984
rect 42061 40987 42119 40993
rect 40828 40944 40834 40956
rect 42061 40953 42073 40987
rect 42107 40953 42119 40987
rect 42061 40947 42119 40953
rect 42334 40944 42340 40996
rect 42392 40984 42398 40996
rect 42720 40984 42748 41083
rect 42904 41052 42932 41083
rect 43162 41080 43168 41083
rect 43220 41120 43226 41132
rect 43898 41120 43904 41132
rect 43220 41092 43267 41120
rect 43859 41092 43904 41120
rect 43220 41080 43226 41092
rect 43898 41080 43904 41092
rect 43956 41080 43962 41132
rect 46569 41123 46627 41129
rect 46569 41089 46581 41123
rect 46615 41120 46627 41123
rect 46658 41120 46664 41132
rect 46615 41092 46664 41120
rect 46615 41089 46627 41092
rect 46569 41083 46627 41089
rect 46658 41080 46664 41092
rect 46716 41080 46722 41132
rect 48314 41080 48320 41132
rect 48372 41120 48378 41132
rect 48501 41123 48559 41129
rect 48501 41120 48513 41123
rect 48372 41092 48513 41120
rect 48372 41080 48378 41092
rect 48501 41089 48513 41092
rect 48547 41089 48559 41123
rect 48501 41083 48559 41089
rect 48705 41092 49281 41120
rect 42978 41052 42984 41064
rect 42904 41024 42984 41052
rect 42978 41012 42984 41024
rect 43036 41012 43042 41064
rect 43809 41055 43867 41061
rect 43809 41021 43821 41055
rect 43855 41021 43867 41055
rect 43809 41015 43867 41021
rect 44269 41055 44327 41061
rect 44269 41021 44281 41055
rect 44315 41052 44327 41055
rect 46293 41055 46351 41061
rect 46293 41052 46305 41055
rect 44315 41024 46305 41052
rect 44315 41021 44327 41024
rect 44269 41015 44327 41021
rect 46293 41021 46305 41024
rect 46339 41021 46351 41055
rect 48705 41052 48733 41092
rect 46293 41015 46351 41021
rect 46492 41024 48733 41052
rect 48777 41055 48835 41061
rect 42392 40956 42748 40984
rect 43257 40987 43315 40993
rect 42392 40944 42398 40956
rect 43257 40953 43269 40987
rect 43303 40984 43315 40987
rect 43824 40984 43852 41015
rect 43303 40956 43852 40984
rect 43303 40953 43315 40956
rect 43257 40947 43315 40953
rect 36630 40876 36636 40928
rect 36688 40916 36694 40928
rect 37550 40916 37556 40928
rect 36688 40888 37556 40916
rect 36688 40876 36694 40888
rect 37550 40876 37556 40888
rect 37608 40876 37614 40928
rect 38102 40876 38108 40928
rect 38160 40916 38166 40928
rect 39301 40919 39359 40925
rect 39301 40916 39313 40919
rect 38160 40888 39313 40916
rect 38160 40876 38166 40888
rect 39301 40885 39313 40888
rect 39347 40885 39359 40919
rect 39301 40879 39359 40885
rect 39666 40876 39672 40928
rect 39724 40916 39730 40928
rect 39945 40919 40003 40925
rect 39945 40916 39957 40919
rect 39724 40888 39957 40916
rect 39724 40876 39730 40888
rect 39945 40885 39957 40888
rect 39991 40885 40003 40919
rect 39945 40879 40003 40885
rect 40037 40919 40095 40925
rect 40037 40885 40049 40919
rect 40083 40916 40095 40919
rect 40126 40916 40132 40928
rect 40083 40888 40132 40916
rect 40083 40885 40095 40888
rect 40037 40879 40095 40885
rect 40126 40876 40132 40888
rect 40184 40876 40190 40928
rect 42242 40876 42248 40928
rect 42300 40916 42306 40928
rect 46492 40916 46520 41024
rect 48777 41021 48789 41055
rect 48823 41052 48835 41055
rect 48866 41052 48872 41064
rect 48823 41024 48872 41052
rect 48823 41021 48835 41024
rect 48777 41015 48835 41021
rect 48866 41012 48872 41024
rect 48924 41012 48930 41064
rect 49253 41052 49281 41092
rect 49326 41080 49332 41132
rect 49384 41120 49390 41132
rect 49602 41120 49608 41132
rect 49384 41092 49608 41120
rect 49384 41080 49390 41092
rect 49602 41080 49608 41092
rect 49660 41080 49666 41132
rect 50246 41052 50252 41064
rect 49253 41024 50252 41052
rect 50246 41012 50252 41024
rect 50304 41012 50310 41064
rect 48406 40944 48412 40996
rect 48464 40984 48470 40996
rect 48593 40987 48651 40993
rect 48593 40984 48605 40987
rect 48464 40956 48605 40984
rect 48464 40944 48470 40956
rect 48593 40953 48605 40956
rect 48639 40984 48651 40987
rect 49602 40984 49608 40996
rect 48639 40956 49608 40984
rect 48639 40953 48651 40956
rect 48593 40947 48651 40953
rect 49602 40944 49608 40956
rect 49660 40944 49666 40996
rect 50724 40984 50752 41160
rect 51718 41148 51724 41200
rect 51776 41188 51782 41200
rect 51776 41160 51821 41188
rect 51776 41148 51782 41160
rect 51902 41148 51908 41200
rect 51960 41188 51966 41200
rect 53009 41191 53067 41197
rect 53009 41188 53021 41191
rect 51960 41160 53021 41188
rect 51960 41148 51966 41160
rect 53009 41157 53021 41160
rect 53055 41188 53067 41191
rect 54386 41188 54392 41200
rect 53055 41160 54392 41188
rect 53055 41157 53067 41160
rect 53009 41151 53067 41157
rect 54386 41148 54392 41160
rect 54444 41188 54450 41200
rect 54754 41188 54760 41200
rect 54444 41160 54760 41188
rect 54444 41148 54450 41160
rect 54754 41148 54760 41160
rect 54812 41148 54818 41200
rect 50798 41080 50804 41132
rect 50856 41120 50862 41132
rect 51077 41123 51135 41129
rect 50856 41092 50901 41120
rect 50856 41080 50862 41092
rect 51077 41089 51089 41123
rect 51123 41120 51135 41123
rect 51537 41123 51595 41129
rect 51537 41120 51549 41123
rect 51123 41092 51549 41120
rect 51123 41089 51135 41092
rect 51077 41083 51135 41089
rect 51537 41089 51549 41092
rect 51583 41120 51595 41123
rect 51626 41120 51632 41132
rect 51583 41092 51632 41120
rect 51583 41089 51595 41092
rect 51537 41083 51595 41089
rect 51626 41080 51632 41092
rect 51684 41080 51690 41132
rect 51810 41129 51816 41132
rect 51809 41083 51816 41129
rect 51868 41120 51874 41132
rect 51868 41092 51909 41120
rect 51810 41080 51816 41083
rect 51868 41080 51874 41092
rect 51994 41080 52000 41132
rect 52052 41120 52058 41132
rect 52273 41123 52331 41129
rect 52273 41120 52285 41123
rect 52052 41092 52285 41120
rect 52052 41080 52058 41092
rect 52273 41089 52285 41092
rect 52319 41120 52331 41123
rect 52362 41120 52368 41132
rect 52319 41092 52368 41120
rect 52319 41089 52331 41092
rect 52273 41083 52331 41089
rect 52362 41080 52368 41092
rect 52420 41080 52426 41132
rect 53834 41120 53840 41132
rect 53747 41092 53840 41120
rect 53834 41080 53840 41092
rect 53892 41120 53898 41132
rect 54018 41120 54024 41132
rect 53892 41092 54024 41120
rect 53892 41080 53898 41092
rect 54018 41080 54024 41092
rect 54076 41080 54082 41132
rect 55232 41129 55260 41228
rect 55585 41225 55597 41259
rect 55631 41256 55643 41259
rect 56226 41256 56232 41268
rect 55631 41228 56232 41256
rect 55631 41225 55643 41228
rect 55585 41219 55643 41225
rect 56226 41216 56232 41228
rect 56284 41216 56290 41268
rect 55217 41123 55275 41129
rect 54409 41092 55168 41120
rect 54409 41052 54437 41092
rect 52656 41024 54437 41052
rect 52656 40984 52684 41024
rect 54478 41012 54484 41064
rect 54536 41052 54542 41064
rect 54662 41052 54668 41064
rect 54536 41024 54668 41052
rect 54536 41012 54542 41024
rect 54662 41012 54668 41024
rect 54720 41012 54726 41064
rect 55140 41061 55168 41092
rect 55217 41089 55229 41123
rect 55263 41089 55275 41123
rect 55217 41083 55275 41089
rect 55125 41055 55183 41061
rect 55125 41021 55137 41055
rect 55171 41052 55183 41055
rect 55582 41052 55588 41064
rect 55171 41024 55588 41052
rect 55171 41021 55183 41024
rect 55125 41015 55183 41021
rect 55582 41012 55588 41024
rect 55640 41012 55646 41064
rect 54570 40984 54576 40996
rect 50724 40956 52684 40984
rect 53116 40956 54576 40984
rect 53116 40928 53144 40956
rect 54570 40944 54576 40956
rect 54628 40944 54634 40996
rect 42300 40888 46520 40916
rect 48685 40919 48743 40925
rect 42300 40876 42306 40888
rect 48685 40885 48697 40919
rect 48731 40916 48743 40919
rect 48958 40916 48964 40928
rect 48731 40888 48964 40916
rect 48731 40885 48743 40888
rect 48685 40879 48743 40885
rect 48958 40876 48964 40888
rect 49016 40876 49022 40928
rect 51077 40919 51135 40925
rect 51077 40885 51089 40919
rect 51123 40916 51135 40919
rect 51166 40916 51172 40928
rect 51123 40888 51172 40916
rect 51123 40885 51135 40888
rect 51077 40879 51135 40885
rect 51166 40876 51172 40888
rect 51224 40876 51230 40928
rect 51537 40919 51595 40925
rect 51537 40885 51549 40919
rect 51583 40916 51595 40919
rect 51994 40916 52000 40928
rect 51583 40888 52000 40916
rect 51583 40885 51595 40888
rect 51537 40879 51595 40885
rect 51994 40876 52000 40888
rect 52052 40876 52058 40928
rect 53098 40916 53104 40928
rect 53059 40888 53104 40916
rect 53098 40876 53104 40888
rect 53156 40876 53162 40928
rect 53926 40876 53932 40928
rect 53984 40916 53990 40928
rect 54021 40919 54079 40925
rect 54021 40916 54033 40919
rect 53984 40888 54033 40916
rect 53984 40876 53990 40888
rect 54021 40885 54033 40888
rect 54067 40885 54079 40919
rect 54021 40879 54079 40885
rect 55030 40876 55036 40928
rect 55088 40916 55094 40928
rect 56045 40919 56103 40925
rect 56045 40916 56057 40919
rect 55088 40888 56057 40916
rect 55088 40876 55094 40888
rect 56045 40885 56057 40888
rect 56091 40916 56103 40919
rect 56597 40919 56655 40925
rect 56597 40916 56609 40919
rect 56091 40888 56609 40916
rect 56091 40885 56103 40888
rect 56045 40879 56103 40885
rect 56597 40885 56609 40888
rect 56643 40885 56655 40919
rect 56597 40879 56655 40885
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 29086 40712 29092 40724
rect 29047 40684 29092 40712
rect 29086 40672 29092 40684
rect 29144 40672 29150 40724
rect 30834 40672 30840 40724
rect 30892 40712 30898 40724
rect 31205 40715 31263 40721
rect 31205 40712 31217 40715
rect 30892 40684 31217 40712
rect 30892 40672 30898 40684
rect 31205 40681 31217 40684
rect 31251 40681 31263 40715
rect 31205 40675 31263 40681
rect 32309 40715 32367 40721
rect 32309 40681 32321 40715
rect 32355 40712 32367 40715
rect 32398 40712 32404 40724
rect 32355 40684 32404 40712
rect 32355 40681 32367 40684
rect 32309 40675 32367 40681
rect 32398 40672 32404 40684
rect 32456 40672 32462 40724
rect 34698 40672 34704 40724
rect 34756 40712 34762 40724
rect 35161 40715 35219 40721
rect 35161 40712 35173 40715
rect 34756 40684 35173 40712
rect 34756 40672 34762 40684
rect 35161 40681 35173 40684
rect 35207 40681 35219 40715
rect 35161 40675 35219 40681
rect 35253 40715 35311 40721
rect 35253 40681 35265 40715
rect 35299 40712 35311 40715
rect 35894 40712 35900 40724
rect 35299 40684 35900 40712
rect 35299 40681 35311 40684
rect 35253 40675 35311 40681
rect 35894 40672 35900 40684
rect 35952 40672 35958 40724
rect 36265 40715 36323 40721
rect 36265 40681 36277 40715
rect 36311 40712 36323 40715
rect 36630 40712 36636 40724
rect 36311 40684 36636 40712
rect 36311 40681 36323 40684
rect 36265 40675 36323 40681
rect 36630 40672 36636 40684
rect 36688 40672 36694 40724
rect 36722 40672 36728 40724
rect 36780 40712 36786 40724
rect 36909 40715 36967 40721
rect 36909 40712 36921 40715
rect 36780 40684 36921 40712
rect 36780 40672 36786 40684
rect 36909 40681 36921 40684
rect 36955 40681 36967 40715
rect 37918 40712 37924 40724
rect 37879 40684 37924 40712
rect 36909 40675 36967 40681
rect 37918 40672 37924 40684
rect 37976 40672 37982 40724
rect 38470 40672 38476 40724
rect 38528 40712 38534 40724
rect 38657 40715 38715 40721
rect 38657 40712 38669 40715
rect 38528 40684 38669 40712
rect 38528 40672 38534 40684
rect 38657 40681 38669 40684
rect 38703 40712 38715 40715
rect 40034 40712 40040 40724
rect 38703 40684 40040 40712
rect 38703 40681 38715 40684
rect 38657 40675 38715 40681
rect 40034 40672 40040 40684
rect 40092 40712 40098 40724
rect 40129 40715 40187 40721
rect 40129 40712 40141 40715
rect 40092 40684 40141 40712
rect 40092 40672 40098 40684
rect 40129 40681 40141 40684
rect 40175 40712 40187 40715
rect 45002 40712 45008 40724
rect 40175 40684 45008 40712
rect 40175 40681 40187 40684
rect 40129 40675 40187 40681
rect 45002 40672 45008 40684
rect 45060 40672 45066 40724
rect 53377 40715 53435 40721
rect 45112 40684 46796 40712
rect 30760 40616 35112 40644
rect 28721 40579 28779 40585
rect 28721 40545 28733 40579
rect 28767 40576 28779 40579
rect 29822 40576 29828 40588
rect 28767 40548 29828 40576
rect 28767 40545 28779 40548
rect 28721 40539 28779 40545
rect 29822 40536 29828 40548
rect 29880 40536 29886 40588
rect 28813 40511 28871 40517
rect 28813 40477 28825 40511
rect 28859 40508 28871 40511
rect 28902 40508 28908 40520
rect 28859 40480 28908 40508
rect 28859 40477 28871 40480
rect 28813 40471 28871 40477
rect 28902 40468 28908 40480
rect 28960 40468 28966 40520
rect 30558 40508 30564 40520
rect 30519 40480 30564 40508
rect 30558 40468 30564 40480
rect 30616 40468 30622 40520
rect 30654 40511 30712 40517
rect 30654 40477 30666 40511
rect 30700 40508 30712 40511
rect 30760 40508 30788 40616
rect 32398 40536 32404 40588
rect 32456 40576 32462 40588
rect 32953 40579 33011 40585
rect 32953 40576 32965 40579
rect 32456 40548 32965 40576
rect 32456 40536 32462 40548
rect 32953 40545 32965 40548
rect 32999 40545 33011 40579
rect 32953 40539 33011 40545
rect 30700 40480 30788 40508
rect 31067 40511 31125 40517
rect 30700 40477 30712 40480
rect 30654 40471 30712 40477
rect 31067 40477 31079 40511
rect 31113 40508 31125 40511
rect 31754 40508 31760 40520
rect 31113 40480 31760 40508
rect 31113 40477 31125 40480
rect 31067 40471 31125 40477
rect 30374 40400 30380 40452
rect 30432 40440 30438 40452
rect 30668 40440 30696 40471
rect 31754 40468 31760 40480
rect 31812 40468 31818 40520
rect 32493 40511 32551 40517
rect 32493 40477 32505 40511
rect 32539 40508 32551 40511
rect 32766 40508 32772 40520
rect 32539 40480 32772 40508
rect 32539 40477 32551 40480
rect 32493 40471 32551 40477
rect 32766 40468 32772 40480
rect 32824 40468 32830 40520
rect 33137 40511 33195 40517
rect 33137 40477 33149 40511
rect 33183 40477 33195 40511
rect 33137 40471 33195 40477
rect 30834 40440 30840 40452
rect 30432 40412 30696 40440
rect 30795 40412 30840 40440
rect 30432 40400 30438 40412
rect 30834 40400 30840 40412
rect 30892 40400 30898 40452
rect 30926 40400 30932 40452
rect 30984 40440 30990 40452
rect 31846 40440 31852 40452
rect 30984 40412 31852 40440
rect 30984 40400 30990 40412
rect 31846 40400 31852 40412
rect 31904 40400 31910 40452
rect 32582 40400 32588 40452
rect 32640 40440 32646 40452
rect 33152 40440 33180 40471
rect 33226 40468 33232 40520
rect 33284 40508 33290 40520
rect 35084 40517 35112 40616
rect 35526 40604 35532 40656
rect 35584 40644 35590 40656
rect 40770 40644 40776 40656
rect 35584 40616 40776 40644
rect 35584 40604 35590 40616
rect 40770 40604 40776 40616
rect 40828 40604 40834 40656
rect 42613 40647 42671 40653
rect 42613 40613 42625 40647
rect 42659 40644 42671 40647
rect 42702 40644 42708 40656
rect 42659 40616 42708 40644
rect 42659 40613 42671 40616
rect 42613 40607 42671 40613
rect 42702 40604 42708 40616
rect 42760 40604 42766 40656
rect 35342 40576 35348 40588
rect 35303 40548 35348 40576
rect 35342 40536 35348 40548
rect 35400 40536 35406 40588
rect 35069 40511 35127 40517
rect 33284 40480 33329 40508
rect 33284 40468 33290 40480
rect 35069 40477 35081 40511
rect 35115 40508 35127 40511
rect 35250 40508 35256 40520
rect 35115 40480 35256 40508
rect 35115 40477 35127 40480
rect 35069 40471 35127 40477
rect 35250 40468 35256 40480
rect 35308 40508 35314 40520
rect 35544 40508 35572 40604
rect 37093 40579 37151 40585
rect 37093 40545 37105 40579
rect 37139 40576 37151 40579
rect 37182 40576 37188 40588
rect 37139 40548 37188 40576
rect 37139 40545 37151 40548
rect 37093 40539 37151 40545
rect 37182 40536 37188 40548
rect 37240 40536 37246 40588
rect 37826 40576 37832 40588
rect 37787 40548 37832 40576
rect 37826 40536 37832 40548
rect 37884 40536 37890 40588
rect 45112 40576 45140 40684
rect 45741 40647 45799 40653
rect 45741 40613 45753 40647
rect 45787 40613 45799 40647
rect 46768 40644 46796 40684
rect 53377 40681 53389 40715
rect 53423 40712 53435 40715
rect 54110 40712 54116 40724
rect 53423 40684 54116 40712
rect 53423 40681 53435 40684
rect 53377 40675 53435 40681
rect 54110 40672 54116 40684
rect 54168 40672 54174 40724
rect 48130 40644 48136 40656
rect 46768 40616 48136 40644
rect 45741 40607 45799 40613
rect 45278 40576 45284 40588
rect 41386 40548 45140 40576
rect 45239 40548 45284 40576
rect 35308 40480 35572 40508
rect 35308 40468 35314 40480
rect 36722 40468 36728 40520
rect 36780 40508 36786 40520
rect 36817 40511 36875 40517
rect 36817 40508 36829 40511
rect 36780 40480 36829 40508
rect 36780 40468 36786 40480
rect 36817 40477 36829 40480
rect 36863 40477 36875 40511
rect 36817 40471 36875 40477
rect 36998 40468 37004 40520
rect 37056 40508 37062 40520
rect 38013 40511 38071 40517
rect 38013 40508 38025 40511
rect 37056 40480 38025 40508
rect 37056 40468 37062 40480
rect 38013 40477 38025 40480
rect 38059 40477 38071 40511
rect 38013 40471 38071 40477
rect 38105 40511 38163 40517
rect 38105 40477 38117 40511
rect 38151 40508 38163 40511
rect 39206 40508 39212 40520
rect 38151 40480 39212 40508
rect 38151 40477 38163 40480
rect 38105 40471 38163 40477
rect 39206 40468 39212 40480
rect 39264 40468 39270 40520
rect 40678 40508 40684 40520
rect 40639 40480 40684 40508
rect 40678 40468 40684 40480
rect 40736 40468 40742 40520
rect 37016 40440 37044 40468
rect 32640 40412 37044 40440
rect 32640 40400 32646 40412
rect 37642 40400 37648 40452
rect 37700 40440 37706 40452
rect 37918 40440 37924 40452
rect 37700 40412 37924 40440
rect 37700 40400 37706 40412
rect 37918 40400 37924 40412
rect 37976 40400 37982 40452
rect 39482 40440 39488 40452
rect 38626 40412 39488 40440
rect 32950 40372 32956 40384
rect 32911 40344 32956 40372
rect 32950 40332 32956 40344
rect 33008 40332 33014 40384
rect 37090 40372 37096 40384
rect 37051 40344 37096 40372
rect 37090 40332 37096 40344
rect 37148 40332 37154 40384
rect 37182 40332 37188 40384
rect 37240 40372 37246 40384
rect 38626 40372 38654 40412
rect 39482 40400 39488 40412
rect 39540 40400 39546 40452
rect 37240 40344 38654 40372
rect 39209 40375 39267 40381
rect 37240 40332 37246 40344
rect 39209 40341 39221 40375
rect 39255 40372 39267 40375
rect 40034 40372 40040 40384
rect 39255 40344 40040 40372
rect 39255 40341 39267 40344
rect 39209 40335 39267 40341
rect 40034 40332 40040 40344
rect 40092 40332 40098 40384
rect 40494 40332 40500 40384
rect 40552 40372 40558 40384
rect 40773 40375 40831 40381
rect 40773 40372 40785 40375
rect 40552 40344 40785 40372
rect 40552 40332 40558 40344
rect 40773 40341 40785 40344
rect 40819 40372 40831 40375
rect 41386 40372 41414 40548
rect 45278 40536 45284 40548
rect 45336 40536 45342 40588
rect 45756 40576 45784 40607
rect 48130 40604 48136 40616
rect 48188 40604 48194 40656
rect 48406 40604 48412 40656
rect 48464 40644 48470 40656
rect 51534 40644 51540 40656
rect 48464 40616 51540 40644
rect 48464 40604 48470 40616
rect 51534 40604 51540 40616
rect 51592 40604 51598 40656
rect 52641 40647 52699 40653
rect 52641 40613 52653 40647
rect 52687 40644 52699 40647
rect 52687 40616 55720 40644
rect 52687 40613 52699 40616
rect 52641 40607 52699 40613
rect 46569 40579 46627 40585
rect 46569 40576 46581 40579
rect 45756 40548 46581 40576
rect 46569 40545 46581 40548
rect 46615 40545 46627 40579
rect 46569 40539 46627 40545
rect 48314 40536 48320 40588
rect 48372 40576 48378 40588
rect 50890 40576 50896 40588
rect 48372 40548 48636 40576
rect 50851 40548 50896 40576
rect 48372 40536 48378 40548
rect 41690 40468 41696 40520
rect 41748 40508 41754 40520
rect 42337 40511 42395 40517
rect 42337 40508 42349 40511
rect 41748 40480 42349 40508
rect 41748 40468 41754 40480
rect 42337 40477 42349 40480
rect 42383 40477 42395 40511
rect 42337 40471 42395 40477
rect 45373 40511 45431 40517
rect 45373 40477 45385 40511
rect 45419 40508 45431 40511
rect 45462 40508 45468 40520
rect 45419 40480 45468 40508
rect 45419 40477 45431 40480
rect 45373 40471 45431 40477
rect 45462 40468 45468 40480
rect 45520 40468 45526 40520
rect 46658 40508 46664 40520
rect 46619 40480 46664 40508
rect 46658 40468 46664 40480
rect 46716 40468 46722 40520
rect 48608 40517 48636 40548
rect 50890 40536 50896 40548
rect 50948 40536 50954 40588
rect 51166 40536 51172 40588
rect 51224 40576 51230 40588
rect 53469 40579 53527 40585
rect 51224 40548 52684 40576
rect 51224 40536 51230 40548
rect 48496 40511 48554 40517
rect 48496 40477 48508 40511
rect 48542 40477 48554 40511
rect 48496 40471 48554 40477
rect 48593 40511 48651 40517
rect 48593 40477 48605 40511
rect 48639 40477 48651 40511
rect 48593 40471 48651 40477
rect 41966 40400 41972 40452
rect 42024 40440 42030 40452
rect 42613 40443 42671 40449
rect 42613 40440 42625 40443
rect 42024 40412 42625 40440
rect 42024 40400 42030 40412
rect 42613 40409 42625 40412
rect 42659 40440 42671 40443
rect 45186 40440 45192 40452
rect 42659 40412 45192 40440
rect 42659 40409 42671 40412
rect 42613 40403 42671 40409
rect 45186 40400 45192 40412
rect 45244 40400 45250 40452
rect 40819 40344 41414 40372
rect 40819 40341 40831 40344
rect 40773 40335 40831 40341
rect 42058 40332 42064 40384
rect 42116 40372 42122 40384
rect 42429 40375 42487 40381
rect 42429 40372 42441 40375
rect 42116 40344 42441 40372
rect 42116 40332 42122 40344
rect 42429 40341 42441 40344
rect 42475 40341 42487 40375
rect 47486 40372 47492 40384
rect 47447 40344 47492 40372
rect 42429 40335 42487 40341
rect 47486 40332 47492 40344
rect 47544 40332 47550 40384
rect 48314 40372 48320 40384
rect 48275 40344 48320 40372
rect 48314 40332 48320 40344
rect 48372 40332 48378 40384
rect 48521 40372 48549 40471
rect 48774 40468 48780 40520
rect 48832 40517 48838 40520
rect 48832 40511 48871 40517
rect 48859 40477 48871 40511
rect 48832 40471 48871 40477
rect 48832 40468 48838 40471
rect 48958 40468 48964 40520
rect 49016 40508 49022 40520
rect 49016 40480 49061 40508
rect 49016 40468 49022 40480
rect 49510 40468 49516 40520
rect 49568 40508 49574 40520
rect 50617 40511 50675 40517
rect 50617 40508 50629 40511
rect 49568 40480 50629 40508
rect 49568 40468 49574 40480
rect 50617 40477 50629 40480
rect 50663 40477 50675 40511
rect 51994 40508 52000 40520
rect 51955 40480 52000 40508
rect 50617 40471 50675 40477
rect 51994 40468 52000 40480
rect 52052 40468 52058 40520
rect 52086 40468 52092 40520
rect 52144 40508 52150 40520
rect 52362 40508 52368 40520
rect 52144 40480 52189 40508
rect 52323 40480 52368 40508
rect 52144 40468 52150 40480
rect 52362 40468 52368 40480
rect 52420 40468 52426 40520
rect 52462 40511 52520 40517
rect 52462 40477 52474 40511
rect 52508 40477 52520 40511
rect 52656 40508 52684 40548
rect 53469 40545 53481 40579
rect 53515 40576 53527 40579
rect 53650 40576 53656 40588
rect 53515 40548 53656 40576
rect 53515 40545 53527 40548
rect 53469 40539 53527 40545
rect 53650 40536 53656 40548
rect 53708 40536 53714 40588
rect 53834 40536 53840 40588
rect 53892 40576 53898 40588
rect 54294 40576 54300 40588
rect 53892 40548 54300 40576
rect 53892 40536 53898 40548
rect 53193 40511 53251 40517
rect 53193 40508 53205 40511
rect 52656 40480 53205 40508
rect 52462 40471 52520 40477
rect 53193 40477 53205 40480
rect 53239 40477 53251 40511
rect 53193 40471 53251 40477
rect 53285 40511 53343 40517
rect 53285 40477 53297 40511
rect 53331 40508 53343 40511
rect 53374 40508 53380 40520
rect 53331 40480 53380 40508
rect 53331 40477 53343 40480
rect 53285 40471 53343 40477
rect 48685 40443 48743 40449
rect 48685 40409 48697 40443
rect 48731 40440 48743 40443
rect 49418 40440 49424 40452
rect 48731 40412 49424 40440
rect 48731 40409 48743 40412
rect 48685 40403 48743 40409
rect 49418 40400 49424 40412
rect 49476 40400 49482 40452
rect 49878 40440 49884 40452
rect 49528 40412 49884 40440
rect 49528 40372 49556 40412
rect 49878 40400 49884 40412
rect 49936 40440 49942 40452
rect 51258 40440 51264 40452
rect 49936 40412 51264 40440
rect 49936 40400 49942 40412
rect 51258 40400 51264 40412
rect 51316 40440 51322 40452
rect 52270 40440 52276 40452
rect 51316 40412 52133 40440
rect 52231 40412 52276 40440
rect 51316 40400 51322 40412
rect 49694 40372 49700 40384
rect 48521 40344 49556 40372
rect 49655 40344 49700 40372
rect 49694 40332 49700 40344
rect 49752 40372 49758 40384
rect 51166 40372 51172 40384
rect 49752 40344 51172 40372
rect 49752 40332 49758 40344
rect 51166 40332 51172 40344
rect 51224 40332 51230 40384
rect 51442 40372 51448 40384
rect 51403 40344 51448 40372
rect 51442 40332 51448 40344
rect 51500 40332 51506 40384
rect 52105 40372 52133 40412
rect 52270 40400 52276 40412
rect 52328 40400 52334 40452
rect 52477 40440 52505 40471
rect 52822 40440 52828 40452
rect 52477 40412 52828 40440
rect 52822 40400 52828 40412
rect 52880 40400 52886 40452
rect 53208 40440 53236 40471
rect 53374 40468 53380 40480
rect 53432 40468 53438 40520
rect 53926 40508 53932 40520
rect 53887 40480 53932 40508
rect 53926 40468 53932 40480
rect 53984 40468 53990 40520
rect 54018 40468 54024 40520
rect 54076 40508 54082 40520
rect 54220 40517 54248 40548
rect 54294 40536 54300 40548
rect 54352 40536 54358 40588
rect 54205 40511 54263 40517
rect 54076 40480 54121 40508
rect 54076 40468 54082 40480
rect 54205 40477 54217 40511
rect 54251 40477 54263 40511
rect 54205 40471 54263 40477
rect 54394 40511 54452 40517
rect 54394 40477 54406 40511
rect 54440 40508 54452 40511
rect 54570 40508 54576 40520
rect 54440 40480 54576 40508
rect 54440 40477 54452 40480
rect 54394 40471 54452 40477
rect 54570 40468 54576 40480
rect 54628 40468 54634 40520
rect 55582 40508 55588 40520
rect 55543 40480 55588 40508
rect 55582 40468 55588 40480
rect 55640 40468 55646 40520
rect 55692 40494 55720 40616
rect 57238 40508 57244 40520
rect 57199 40480 57244 40508
rect 57238 40468 57244 40480
rect 57296 40468 57302 40520
rect 57422 40508 57428 40520
rect 57383 40480 57428 40508
rect 57422 40468 57428 40480
rect 57480 40468 57486 40520
rect 54036 40440 54064 40468
rect 53208 40412 54064 40440
rect 54297 40443 54355 40449
rect 54297 40409 54309 40443
rect 54343 40440 54355 40443
rect 54478 40440 54484 40452
rect 54343 40412 54484 40440
rect 54343 40409 54355 40412
rect 54297 40403 54355 40409
rect 54478 40400 54484 40412
rect 54536 40440 54542 40452
rect 55030 40440 55036 40452
rect 54536 40412 55036 40440
rect 54536 40400 54542 40412
rect 55030 40400 55036 40412
rect 55088 40400 55094 40452
rect 56594 40440 56600 40452
rect 56555 40412 56600 40440
rect 56594 40400 56600 40412
rect 56652 40400 56658 40452
rect 53098 40372 53104 40384
rect 52105 40344 53104 40372
rect 53098 40332 53104 40344
rect 53156 40332 53162 40384
rect 54573 40375 54631 40381
rect 54573 40341 54585 40375
rect 54619 40372 54631 40375
rect 54846 40372 54852 40384
rect 54619 40344 54852 40372
rect 54619 40341 54631 40344
rect 54573 40335 54631 40341
rect 54846 40332 54852 40344
rect 54904 40332 54910 40384
rect 58250 40372 58256 40384
rect 58211 40344 58256 40372
rect 58250 40332 58256 40344
rect 58308 40332 58314 40384
rect 1104 40282 58880 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 35594 40282
rect 35646 40230 35658 40282
rect 35710 40230 35722 40282
rect 35774 40230 35786 40282
rect 35838 40230 35850 40282
rect 35902 40230 58880 40282
rect 1104 40208 58880 40230
rect 30834 40128 30840 40180
rect 30892 40168 30898 40180
rect 31570 40168 31576 40180
rect 30892 40140 31576 40168
rect 30892 40128 30898 40140
rect 31036 40109 31064 40140
rect 31570 40128 31576 40140
rect 31628 40168 31634 40180
rect 31628 40140 32720 40168
rect 31628 40128 31634 40140
rect 30285 40103 30343 40109
rect 30285 40069 30297 40103
rect 30331 40100 30343 40103
rect 31021 40103 31079 40109
rect 30331 40072 30788 40100
rect 30331 40069 30343 40072
rect 30285 40063 30343 40069
rect 30009 40035 30067 40041
rect 30009 40001 30021 40035
rect 30055 40032 30067 40035
rect 30650 40032 30656 40044
rect 30055 40004 30656 40032
rect 30055 40001 30067 40004
rect 30009 39995 30067 40001
rect 30650 39992 30656 40004
rect 30708 39992 30714 40044
rect 30760 40041 30788 40072
rect 31021 40069 31033 40103
rect 31067 40069 31079 40103
rect 31754 40100 31760 40112
rect 31021 40063 31079 40069
rect 31404 40072 31760 40100
rect 30926 40041 30932 40044
rect 30745 40035 30803 40041
rect 30745 40001 30757 40035
rect 30791 40001 30803 40035
rect 30745 39995 30803 40001
rect 30893 40035 30932 40041
rect 30893 40001 30905 40035
rect 30893 39995 30932 40001
rect 30926 39992 30932 39995
rect 30984 39992 30990 40044
rect 31110 39992 31116 40044
rect 31168 40032 31174 40044
rect 31251 40035 31309 40041
rect 31168 40004 31213 40032
rect 31168 39992 31174 40004
rect 31251 40001 31263 40035
rect 31297 40032 31309 40035
rect 31404 40032 31432 40072
rect 31754 40060 31760 40072
rect 31812 40060 31818 40112
rect 32692 40109 32720 40140
rect 38102 40128 38108 40180
rect 38160 40168 38166 40180
rect 40402 40168 40408 40180
rect 38160 40140 40408 40168
rect 38160 40128 38166 40140
rect 40402 40128 40408 40140
rect 40460 40128 40466 40180
rect 41870 40171 41928 40177
rect 41386 40140 41828 40168
rect 32585 40103 32643 40109
rect 32585 40100 32597 40103
rect 31864 40072 32597 40100
rect 31864 40032 31892 40072
rect 32585 40069 32597 40072
rect 32631 40069 32643 40103
rect 32585 40063 32643 40069
rect 32677 40103 32735 40109
rect 32677 40069 32689 40103
rect 32723 40069 32735 40103
rect 33226 40100 33232 40112
rect 32677 40063 32735 40069
rect 32876 40072 33232 40100
rect 32490 40041 32496 40044
rect 32488 40032 32496 40041
rect 31297 40004 31432 40032
rect 31726 40004 31892 40032
rect 32451 40004 32496 40032
rect 31297 40001 31309 40004
rect 31251 39995 31309 40001
rect 29178 39924 29184 39976
rect 29236 39964 29242 39976
rect 30285 39967 30343 39973
rect 30285 39964 30297 39967
rect 29236 39936 30297 39964
rect 29236 39924 29242 39936
rect 30285 39933 30297 39936
rect 30331 39933 30343 39967
rect 30285 39927 30343 39933
rect 30374 39924 30380 39976
rect 30432 39964 30438 39976
rect 31726 39964 31754 40004
rect 32488 39995 32496 40004
rect 32490 39992 32496 39995
rect 32548 39992 32554 40044
rect 32876 40041 32904 40072
rect 33226 40060 33232 40072
rect 33284 40100 33290 40112
rect 34606 40100 34612 40112
rect 33284 40072 34612 40100
rect 33284 40060 33290 40072
rect 34606 40060 34612 40072
rect 34664 40060 34670 40112
rect 37734 40060 37740 40112
rect 37792 40100 37798 40112
rect 41386 40100 41414 40140
rect 41800 40109 41828 40140
rect 41870 40137 41882 40171
rect 41916 40168 41928 40171
rect 42978 40168 42984 40180
rect 41916 40140 42288 40168
rect 41916 40137 41928 40140
rect 41870 40131 41928 40137
rect 37792 40072 37837 40100
rect 38672 40072 41414 40100
rect 41785 40103 41843 40109
rect 37792 40060 37798 40072
rect 32860 40035 32918 40041
rect 32860 40001 32872 40035
rect 32906 40001 32918 40035
rect 32860 39995 32918 40001
rect 32950 39992 32956 40044
rect 33008 40032 33014 40044
rect 33594 40032 33600 40044
rect 33008 40004 33053 40032
rect 33555 40004 33600 40032
rect 33008 39992 33014 40004
rect 33594 39992 33600 40004
rect 33652 39992 33658 40044
rect 36078 40032 36084 40044
rect 36039 40004 36084 40032
rect 36078 39992 36084 40004
rect 36136 39992 36142 40044
rect 37090 39992 37096 40044
rect 37148 40032 37154 40044
rect 37642 40041 37648 40044
rect 37450 40035 37508 40041
rect 37450 40032 37462 40035
rect 37148 40004 37462 40032
rect 37148 39992 37154 40004
rect 37450 40001 37462 40004
rect 37496 40001 37508 40035
rect 37450 39995 37508 40001
rect 37609 40035 37648 40041
rect 37609 40001 37621 40035
rect 37609 39995 37648 40001
rect 37642 39992 37648 39995
rect 37700 39992 37706 40044
rect 37829 40035 37887 40041
rect 37829 40032 37841 40035
rect 37752 40004 37841 40032
rect 33502 39964 33508 39976
rect 30432 39936 31754 39964
rect 33463 39936 33508 39964
rect 30432 39924 30438 39936
rect 33502 39924 33508 39936
rect 33560 39924 33566 39976
rect 34054 39924 34060 39976
rect 34112 39964 34118 39976
rect 35897 39967 35955 39973
rect 35897 39964 35909 39967
rect 34112 39936 35909 39964
rect 34112 39924 34118 39936
rect 35897 39933 35909 39936
rect 35943 39933 35955 39967
rect 35897 39927 35955 39933
rect 36817 39967 36875 39973
rect 36817 39933 36829 39967
rect 36863 39933 36875 39967
rect 36817 39927 36875 39933
rect 31386 39896 31392 39908
rect 31347 39868 31392 39896
rect 31386 39856 31392 39868
rect 31444 39856 31450 39908
rect 32306 39896 32312 39908
rect 32267 39868 32312 39896
rect 32306 39856 32312 39868
rect 32364 39856 32370 39908
rect 33962 39896 33968 39908
rect 33923 39868 33968 39896
rect 33962 39856 33968 39868
rect 34020 39856 34026 39908
rect 28994 39788 29000 39840
rect 29052 39828 29058 39840
rect 30101 39831 30159 39837
rect 30101 39828 30113 39831
rect 29052 39800 30113 39828
rect 29052 39788 29058 39800
rect 30101 39797 30113 39800
rect 30147 39828 30159 39831
rect 32214 39828 32220 39840
rect 30147 39800 32220 39828
rect 30147 39797 30159 39800
rect 30101 39791 30159 39797
rect 32214 39788 32220 39800
rect 32272 39788 32278 39840
rect 35250 39788 35256 39840
rect 35308 39828 35314 39840
rect 35526 39828 35532 39840
rect 35308 39800 35532 39828
rect 35308 39788 35314 39800
rect 35526 39788 35532 39800
rect 35584 39788 35590 39840
rect 36832 39828 36860 39927
rect 36906 39856 36912 39908
rect 36964 39896 36970 39908
rect 37752 39896 37780 40004
rect 37829 40001 37841 40004
rect 37875 40001 37887 40035
rect 37829 39995 37887 40001
rect 37918 39992 37924 40044
rect 37976 40041 37982 40044
rect 37976 40035 38025 40041
rect 37976 40001 37979 40035
rect 38013 40032 38025 40035
rect 38562 40032 38568 40044
rect 38013 40004 38568 40032
rect 38013 40001 38025 40004
rect 37976 39995 38025 40001
rect 37976 39992 37982 39995
rect 38562 39992 38568 40004
rect 38620 39992 38626 40044
rect 38102 39924 38108 39976
rect 38160 39964 38166 39976
rect 38672 39964 38700 40072
rect 41785 40069 41797 40103
rect 41831 40069 41843 40103
rect 41966 40100 41972 40112
rect 41927 40072 41972 40100
rect 41785 40063 41843 40069
rect 38838 39992 38844 40044
rect 38896 40032 38902 40044
rect 38933 40035 38991 40041
rect 38933 40032 38945 40035
rect 38896 40004 38945 40032
rect 38896 39992 38902 40004
rect 38933 40001 38945 40004
rect 38979 40001 38991 40035
rect 39850 40032 39856 40044
rect 39811 40004 39856 40032
rect 38933 39995 38991 40001
rect 39850 39992 39856 40004
rect 39908 39992 39914 40044
rect 41690 40032 41696 40044
rect 41651 40004 41696 40032
rect 41690 39992 41696 40004
rect 41748 39992 41754 40044
rect 38160 39936 38700 39964
rect 41800 39964 41828 40063
rect 41966 40060 41972 40072
rect 42024 40060 42030 40112
rect 42260 40032 42288 40140
rect 42904 40140 42984 40168
rect 42334 40060 42340 40112
rect 42392 40100 42398 40112
rect 42904 40109 42932 40140
rect 42978 40128 42984 40140
rect 43036 40128 43042 40180
rect 43257 40171 43315 40177
rect 43257 40137 43269 40171
rect 43303 40137 43315 40171
rect 43257 40131 43315 40137
rect 44269 40171 44327 40177
rect 44269 40137 44281 40171
rect 44315 40168 44327 40171
rect 45278 40168 45284 40180
rect 44315 40140 45284 40168
rect 44315 40137 44327 40140
rect 44269 40131 44327 40137
rect 42889 40103 42947 40109
rect 42392 40072 42840 40100
rect 42392 40060 42398 40072
rect 42613 40035 42671 40041
rect 42613 40032 42625 40035
rect 42260 40004 42625 40032
rect 42613 40001 42625 40004
rect 42659 40001 42671 40035
rect 42613 39995 42671 40001
rect 42706 40035 42764 40041
rect 42706 40001 42718 40035
rect 42752 40001 42764 40035
rect 42812 40032 42840 40072
rect 42889 40069 42901 40103
rect 42935 40069 42947 40103
rect 42889 40063 42947 40069
rect 43162 40041 43168 40044
rect 42981 40035 43039 40041
rect 42981 40032 42993 40035
rect 42812 40004 42993 40032
rect 42706 39995 42764 40001
rect 42981 40001 42993 40004
rect 43027 40001 43039 40035
rect 42981 39995 43039 40001
rect 43119 40035 43168 40041
rect 43119 40001 43131 40035
rect 43165 40001 43168 40035
rect 43119 39995 43168 40001
rect 42518 39964 42524 39976
rect 41800 39936 42524 39964
rect 38160 39924 38166 39936
rect 42518 39924 42524 39936
rect 42576 39964 42582 39976
rect 42720 39964 42748 39995
rect 43162 39992 43168 39995
rect 43220 39992 43226 40044
rect 43272 40032 43300 40131
rect 45278 40128 45284 40140
rect 45336 40128 45342 40180
rect 47486 40128 47492 40180
rect 47544 40168 47550 40180
rect 47544 40140 53880 40168
rect 47544 40128 47550 40140
rect 48314 40060 48320 40112
rect 48372 40100 48378 40112
rect 48372 40072 48636 40100
rect 48372 40060 48378 40072
rect 43901 40035 43959 40041
rect 43901 40032 43913 40035
rect 43272 40004 43913 40032
rect 43901 40001 43913 40004
rect 43947 40001 43959 40035
rect 43901 39995 43959 40001
rect 44450 39992 44456 40044
rect 44508 40032 44514 40044
rect 46753 40035 46811 40041
rect 46753 40032 46765 40035
rect 44508 40004 46765 40032
rect 44508 39992 44514 40004
rect 46753 40001 46765 40004
rect 46799 40032 46811 40035
rect 47026 40032 47032 40044
rect 46799 40004 47032 40032
rect 46799 40001 46811 40004
rect 46753 39995 46811 40001
rect 47026 39992 47032 40004
rect 47084 39992 47090 40044
rect 48608 40041 48636 40072
rect 49510 40060 49516 40112
rect 49568 40100 49574 40112
rect 50985 40103 51043 40109
rect 49568 40072 49648 40100
rect 49568 40060 49574 40072
rect 49620 40041 49648 40072
rect 50985 40069 50997 40103
rect 51031 40100 51043 40103
rect 53374 40100 53380 40112
rect 51031 40072 53380 40100
rect 51031 40069 51043 40072
rect 50985 40063 51043 40069
rect 53374 40060 53380 40072
rect 53432 40060 53438 40112
rect 53558 40060 53564 40112
rect 53616 40100 53622 40112
rect 53852 40100 53880 40140
rect 53926 40128 53932 40180
rect 53984 40168 53990 40180
rect 54021 40171 54079 40177
rect 54021 40168 54033 40171
rect 53984 40140 54033 40168
rect 53984 40128 53990 40140
rect 54021 40137 54033 40140
rect 54067 40137 54079 40171
rect 54021 40131 54079 40137
rect 54110 40128 54116 40180
rect 54168 40168 54174 40180
rect 54662 40168 54668 40180
rect 54168 40140 54668 40168
rect 54168 40128 54174 40140
rect 54662 40128 54668 40140
rect 54720 40128 54726 40180
rect 57149 40171 57207 40177
rect 57149 40137 57161 40171
rect 57195 40168 57207 40171
rect 57238 40168 57244 40180
rect 57195 40140 57244 40168
rect 57195 40137 57207 40140
rect 57149 40131 57207 40137
rect 57238 40128 57244 40140
rect 57296 40128 57302 40180
rect 55674 40100 55680 40112
rect 53616 40072 53788 40100
rect 53852 40072 55680 40100
rect 53616 40060 53622 40072
rect 48593 40035 48651 40041
rect 48593 40001 48605 40035
rect 48639 40001 48651 40035
rect 48593 39995 48651 40001
rect 49605 40035 49663 40041
rect 49605 40001 49617 40035
rect 49651 40001 49663 40035
rect 49605 39995 49663 40001
rect 50246 39992 50252 40044
rect 50304 40032 50310 40044
rect 51905 40035 51963 40041
rect 51905 40032 51917 40035
rect 50304 40004 51917 40032
rect 50304 39992 50310 40004
rect 51905 40001 51917 40004
rect 51951 40032 51963 40035
rect 52086 40032 52092 40044
rect 51951 40004 52092 40032
rect 51951 40001 51963 40004
rect 51905 39995 51963 40001
rect 52086 39992 52092 40004
rect 52144 39992 52150 40044
rect 53009 40035 53067 40041
rect 53009 40001 53021 40035
rect 53055 40032 53067 40035
rect 53650 40032 53656 40044
rect 53055 40004 53656 40032
rect 53055 40001 53067 40004
rect 53009 39995 53067 40001
rect 53650 39992 53656 40004
rect 53708 39992 53714 40044
rect 53760 40041 53788 40072
rect 53745 40035 53803 40041
rect 53745 40001 53757 40035
rect 53791 40032 53803 40035
rect 54110 40032 54116 40044
rect 53791 40004 54116 40032
rect 53791 40001 53803 40004
rect 53745 39995 53803 40001
rect 54110 39992 54116 40004
rect 54168 40032 54174 40044
rect 54478 40032 54484 40044
rect 54168 40004 54484 40032
rect 54168 39992 54174 40004
rect 54478 39992 54484 40004
rect 54536 39992 54542 40044
rect 54956 40041 54984 40072
rect 55674 40060 55680 40072
rect 55732 40060 55738 40112
rect 54941 40035 54999 40041
rect 54941 40001 54953 40035
rect 54987 40001 54999 40035
rect 54941 39995 54999 40001
rect 56594 39992 56600 40044
rect 56652 40032 56658 40044
rect 56781 40035 56839 40041
rect 56781 40032 56793 40035
rect 56652 40004 56793 40032
rect 56652 39992 56658 40004
rect 56781 40001 56793 40004
rect 56827 40032 56839 40035
rect 57238 40032 57244 40044
rect 56827 40004 57244 40032
rect 56827 40001 56839 40004
rect 56781 39995 56839 40001
rect 57238 39992 57244 40004
rect 57296 39992 57302 40044
rect 42576 39936 42748 39964
rect 42576 39924 42582 39936
rect 43530 39924 43536 39976
rect 43588 39964 43594 39976
rect 43809 39967 43867 39973
rect 43809 39964 43821 39967
rect 43588 39936 43821 39964
rect 43588 39924 43594 39936
rect 43809 39933 43821 39936
rect 43855 39933 43867 39967
rect 43809 39927 43867 39933
rect 48314 39924 48320 39976
rect 48372 39964 48378 39976
rect 48501 39967 48559 39973
rect 48501 39964 48513 39967
rect 48372 39936 48513 39964
rect 48372 39924 48378 39936
rect 48501 39933 48513 39936
rect 48547 39933 48559 39967
rect 49513 39967 49571 39973
rect 49513 39964 49525 39967
rect 48501 39927 48559 39933
rect 48976 39936 49525 39964
rect 40773 39899 40831 39905
rect 36964 39868 37780 39896
rect 37982 39868 38654 39896
rect 36964 39856 36970 39868
rect 37982 39828 38010 39868
rect 38102 39828 38108 39840
rect 36832 39800 38010 39828
rect 38063 39800 38108 39828
rect 38102 39788 38108 39800
rect 38160 39788 38166 39840
rect 38626 39828 38654 39868
rect 40773 39865 40785 39899
rect 40819 39896 40831 39899
rect 46658 39896 46664 39908
rect 40819 39868 46664 39896
rect 40819 39865 40831 39868
rect 40773 39859 40831 39865
rect 46658 39856 46664 39868
rect 46716 39856 46722 39908
rect 48976 39905 49004 39936
rect 49513 39933 49525 39936
rect 49559 39933 49571 39967
rect 51261 39967 51319 39973
rect 51261 39964 51273 39967
rect 49513 39927 49571 39933
rect 49620 39936 51273 39964
rect 49620 39908 49648 39936
rect 51261 39933 51273 39936
rect 51307 39964 51319 39967
rect 52914 39964 52920 39976
rect 51307 39936 52920 39964
rect 51307 39933 51319 39936
rect 51261 39927 51319 39933
rect 52914 39924 52920 39936
rect 52972 39924 52978 39976
rect 54021 39967 54079 39973
rect 54021 39964 54033 39967
rect 53576 39936 54033 39964
rect 53576 39908 53604 39936
rect 54021 39933 54033 39936
rect 54067 39933 54079 39967
rect 54846 39964 54852 39976
rect 54807 39936 54852 39964
rect 54021 39927 54079 39933
rect 54846 39924 54852 39936
rect 54904 39924 54910 39976
rect 56689 39967 56747 39973
rect 56689 39964 56701 39967
rect 55324 39936 56701 39964
rect 48961 39899 49019 39905
rect 48961 39865 48973 39899
rect 49007 39865 49019 39899
rect 48961 39859 49019 39865
rect 49602 39856 49608 39908
rect 49660 39856 49666 39908
rect 49973 39899 50031 39905
rect 49973 39865 49985 39899
rect 50019 39896 50031 39899
rect 50154 39896 50160 39908
rect 50019 39868 50160 39896
rect 50019 39865 50031 39868
rect 49973 39859 50031 39865
rect 50154 39856 50160 39868
rect 50212 39856 50218 39908
rect 53190 39896 53196 39908
rect 53103 39868 53196 39896
rect 53190 39856 53196 39868
rect 53248 39896 53254 39908
rect 53558 39896 53564 39908
rect 53248 39868 53564 39896
rect 53248 39856 53254 39868
rect 53558 39856 53564 39868
rect 53616 39856 53622 39908
rect 55324 39905 55352 39936
rect 56689 39933 56701 39936
rect 56735 39933 56747 39967
rect 56689 39927 56747 39933
rect 55309 39899 55367 39905
rect 55309 39865 55321 39899
rect 55355 39865 55367 39899
rect 55309 39859 55367 39865
rect 43898 39828 43904 39840
rect 38626 39800 43904 39828
rect 43898 39788 43904 39800
rect 43956 39788 43962 39840
rect 47670 39788 47676 39840
rect 47728 39828 47734 39840
rect 47765 39831 47823 39837
rect 47765 39828 47777 39831
rect 47728 39800 47777 39828
rect 47728 39788 47734 39800
rect 47765 39797 47777 39800
rect 47811 39828 47823 39831
rect 51718 39828 51724 39840
rect 47811 39800 51724 39828
rect 47811 39797 47823 39800
rect 47765 39791 47823 39797
rect 51718 39788 51724 39800
rect 51776 39788 51782 39840
rect 53374 39788 53380 39840
rect 53432 39828 53438 39840
rect 53837 39831 53895 39837
rect 53837 39828 53849 39831
rect 53432 39800 53849 39828
rect 53432 39788 53438 39800
rect 53837 39797 53849 39800
rect 53883 39797 53895 39831
rect 53837 39791 53895 39797
rect 55582 39788 55588 39840
rect 55640 39828 55646 39840
rect 55769 39831 55827 39837
rect 55769 39828 55781 39831
rect 55640 39800 55781 39828
rect 55640 39788 55646 39800
rect 55769 39797 55781 39800
rect 55815 39797 55827 39831
rect 55769 39791 55827 39797
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 28994 39624 29000 39636
rect 28955 39596 29000 39624
rect 28994 39584 29000 39596
rect 29052 39584 29058 39636
rect 30650 39584 30656 39636
rect 30708 39624 30714 39636
rect 31386 39624 31392 39636
rect 30708 39596 31392 39624
rect 30708 39584 30714 39596
rect 31386 39584 31392 39596
rect 31444 39584 31450 39636
rect 31665 39627 31723 39633
rect 31665 39593 31677 39627
rect 31711 39624 31723 39627
rect 31846 39624 31852 39636
rect 31711 39596 31852 39624
rect 31711 39593 31723 39596
rect 31665 39587 31723 39593
rect 31846 39584 31852 39596
rect 31904 39584 31910 39636
rect 32582 39624 32588 39636
rect 32543 39596 32588 39624
rect 32582 39584 32588 39596
rect 32640 39584 32646 39636
rect 34054 39624 34060 39636
rect 34015 39596 34060 39624
rect 34054 39584 34060 39596
rect 34112 39584 34118 39636
rect 36078 39624 36084 39636
rect 36039 39596 36084 39624
rect 36078 39584 36084 39596
rect 36136 39584 36142 39636
rect 36998 39624 37004 39636
rect 36959 39596 37004 39624
rect 36998 39584 37004 39596
rect 37056 39584 37062 39636
rect 46492 39596 53880 39624
rect 29089 39559 29147 39565
rect 29089 39525 29101 39559
rect 29135 39556 29147 39559
rect 30558 39556 30564 39568
rect 29135 39528 30564 39556
rect 29135 39525 29147 39528
rect 29089 39519 29147 39525
rect 30558 39516 30564 39528
rect 30616 39516 30622 39568
rect 37642 39556 37648 39568
rect 35820 39528 37648 39556
rect 29178 39488 29184 39500
rect 29139 39460 29184 39488
rect 29178 39448 29184 39460
rect 29236 39448 29242 39500
rect 33870 39488 33876 39500
rect 33831 39460 33876 39488
rect 33870 39448 33876 39460
rect 33928 39448 33934 39500
rect 35250 39448 35256 39500
rect 35308 39488 35314 39500
rect 35820 39488 35848 39528
rect 37642 39516 37648 39528
rect 37700 39516 37706 39568
rect 37734 39516 37740 39568
rect 37792 39556 37798 39568
rect 38286 39556 38292 39568
rect 37792 39528 38292 39556
rect 37792 39516 37798 39528
rect 38286 39516 38292 39528
rect 38344 39516 38350 39568
rect 39485 39559 39543 39565
rect 39485 39525 39497 39559
rect 39531 39556 39543 39559
rect 39942 39556 39948 39568
rect 39531 39528 39948 39556
rect 39531 39525 39543 39528
rect 39485 39519 39543 39525
rect 39942 39516 39948 39528
rect 40000 39516 40006 39568
rect 40402 39516 40408 39568
rect 40460 39556 40466 39568
rect 40678 39556 40684 39568
rect 40460 39528 40684 39556
rect 40460 39516 40466 39528
rect 40678 39516 40684 39528
rect 40736 39556 40742 39568
rect 40736 39528 42012 39556
rect 40736 39516 40742 39528
rect 35308 39460 35848 39488
rect 35308 39448 35314 39460
rect 28905 39423 28963 39429
rect 28905 39389 28917 39423
rect 28951 39389 28963 39423
rect 29822 39420 29828 39432
rect 29783 39392 29828 39420
rect 28905 39383 28963 39389
rect 28920 39352 28948 39383
rect 29822 39380 29828 39392
rect 29880 39380 29886 39432
rect 30650 39420 30656 39432
rect 30498 39392 30656 39420
rect 30650 39380 30656 39392
rect 30708 39380 30714 39432
rect 30837 39423 30895 39429
rect 30837 39389 30849 39423
rect 30883 39420 30895 39423
rect 33502 39420 33508 39432
rect 30883 39392 33508 39420
rect 30883 39389 30895 39392
rect 30837 39383 30895 39389
rect 33502 39380 33508 39392
rect 33560 39420 33566 39432
rect 33781 39423 33839 39429
rect 33781 39420 33793 39423
rect 33560 39392 33793 39420
rect 33560 39380 33566 39392
rect 33781 39389 33793 39392
rect 33827 39389 33839 39423
rect 35434 39420 35440 39432
rect 35395 39392 35440 39420
rect 33781 39383 33839 39389
rect 35434 39380 35440 39392
rect 35492 39380 35498 39432
rect 35526 39380 35532 39432
rect 35584 39420 35590 39432
rect 35820 39429 35848 39460
rect 36817 39491 36875 39497
rect 36817 39457 36829 39491
rect 36863 39488 36875 39491
rect 37826 39488 37832 39500
rect 36863 39460 37832 39488
rect 36863 39457 36875 39460
rect 36817 39451 36875 39457
rect 37826 39448 37832 39460
rect 37884 39448 37890 39500
rect 38102 39488 38108 39500
rect 38063 39460 38108 39488
rect 38102 39448 38108 39460
rect 38160 39448 38166 39500
rect 38838 39488 38844 39500
rect 38799 39460 38844 39488
rect 38838 39448 38844 39460
rect 38896 39448 38902 39500
rect 40954 39448 40960 39500
rect 41012 39488 41018 39500
rect 41012 39460 41552 39488
rect 41012 39448 41018 39460
rect 35986 39429 35992 39432
rect 35805 39423 35863 39429
rect 35584 39392 35629 39420
rect 35584 39380 35590 39392
rect 35805 39389 35817 39423
rect 35851 39389 35863 39423
rect 35805 39383 35863 39389
rect 35943 39423 35992 39429
rect 35943 39389 35955 39423
rect 35989 39389 35992 39423
rect 35943 39383 35992 39389
rect 35986 39380 35992 39383
rect 36044 39380 36050 39432
rect 36906 39380 36912 39432
rect 36964 39420 36970 39432
rect 37093 39423 37151 39429
rect 37093 39420 37105 39423
rect 36964 39392 37105 39420
rect 36964 39380 36970 39392
rect 37093 39389 37105 39392
rect 37139 39389 37151 39423
rect 37093 39383 37151 39389
rect 38013 39423 38071 39429
rect 38013 39389 38025 39423
rect 38059 39389 38071 39423
rect 38013 39383 38071 39389
rect 39301 39423 39359 39429
rect 39301 39389 39313 39423
rect 39347 39389 39359 39423
rect 39301 39383 39359 39389
rect 39485 39423 39543 39429
rect 39485 39389 39497 39423
rect 39531 39420 39543 39423
rect 39574 39420 39580 39432
rect 39531 39392 39580 39420
rect 39531 39389 39543 39392
rect 39485 39383 39543 39389
rect 30374 39352 30380 39364
rect 28920 39324 30380 39352
rect 30374 39312 30380 39324
rect 30432 39352 30438 39364
rect 30558 39352 30564 39364
rect 30432 39324 30564 39352
rect 30432 39312 30438 39324
rect 30558 39312 30564 39324
rect 30616 39312 30622 39364
rect 31386 39352 31392 39364
rect 31347 39324 31392 39352
rect 31386 39312 31392 39324
rect 31444 39312 31450 39364
rect 32306 39352 32312 39364
rect 32267 39324 32312 39352
rect 32306 39312 32312 39324
rect 32364 39312 32370 39364
rect 34790 39312 34796 39364
rect 34848 39352 34854 39364
rect 35713 39355 35771 39361
rect 35713 39352 35725 39355
rect 34848 39324 35725 39352
rect 34848 39312 34854 39324
rect 35713 39321 35725 39324
rect 35759 39321 35771 39355
rect 38028 39352 38056 39383
rect 35713 39315 35771 39321
rect 36004 39324 38056 39352
rect 39316 39352 39344 39383
rect 39574 39380 39580 39392
rect 39632 39380 39638 39432
rect 39850 39380 39856 39432
rect 39908 39420 39914 39432
rect 40129 39423 40187 39429
rect 40129 39420 40141 39423
rect 39908 39392 40141 39420
rect 39908 39380 39914 39392
rect 40129 39389 40141 39392
rect 40175 39389 40187 39423
rect 41524 39420 41552 39460
rect 41984 39429 42012 39528
rect 42150 39516 42156 39568
rect 42208 39556 42214 39568
rect 43349 39559 43407 39565
rect 42208 39528 42288 39556
rect 42208 39516 42214 39528
rect 41780 39423 41838 39429
rect 40802 39392 41414 39420
rect 41524 39414 41739 39420
rect 41780 39414 41792 39423
rect 41524 39392 41792 39414
rect 40129 39383 40187 39389
rect 39666 39352 39672 39364
rect 39316 39324 39672 39352
rect 34422 39244 34428 39296
rect 34480 39284 34486 39296
rect 36004 39284 36032 39324
rect 39666 39312 39672 39324
rect 39724 39312 39730 39364
rect 41141 39355 41199 39361
rect 41141 39321 41153 39355
rect 41187 39321 41199 39355
rect 41386 39352 41414 39392
rect 41711 39389 41792 39392
rect 41826 39389 41838 39423
rect 41711 39386 41838 39389
rect 41780 39383 41838 39386
rect 41969 39423 42027 39429
rect 41969 39389 41981 39423
rect 42015 39389 42027 39423
rect 41969 39383 42027 39389
rect 42058 39380 42064 39432
rect 42116 39430 42122 39432
rect 42116 39429 42140 39430
rect 42260 39429 42288 39528
rect 43349 39525 43361 39559
rect 43395 39525 43407 39559
rect 43349 39519 43407 39525
rect 44637 39559 44695 39565
rect 44637 39525 44649 39559
rect 44683 39525 44695 39559
rect 44637 39519 44695 39525
rect 42518 39448 42524 39500
rect 42576 39488 42582 39500
rect 43364 39488 43392 39519
rect 44177 39491 44235 39497
rect 44177 39488 44189 39491
rect 42576 39460 43116 39488
rect 43364 39460 44189 39488
rect 42576 39448 42582 39460
rect 42116 39423 42155 39429
rect 42143 39389 42155 39423
rect 42116 39383 42155 39389
rect 42256 39423 42314 39429
rect 42256 39389 42268 39423
rect 42302 39389 42314 39423
rect 42702 39420 42708 39432
rect 42663 39392 42708 39420
rect 42256 39383 42314 39389
rect 42116 39380 42122 39383
rect 42702 39380 42708 39392
rect 42760 39380 42766 39432
rect 42794 39380 42800 39432
rect 42852 39429 42858 39432
rect 43088 39429 43116 39460
rect 44177 39457 44189 39460
rect 44223 39457 44235 39491
rect 44652 39488 44680 39519
rect 46492 39497 46520 39596
rect 47213 39559 47271 39565
rect 47213 39525 47225 39559
rect 47259 39525 47271 39559
rect 47213 39519 47271 39525
rect 48685 39559 48743 39565
rect 48685 39525 48697 39559
rect 48731 39556 48743 39559
rect 49786 39556 49792 39568
rect 48731 39528 49792 39556
rect 48731 39525 48743 39528
rect 48685 39519 48743 39525
rect 45557 39491 45615 39497
rect 45557 39488 45569 39491
rect 44652 39460 45569 39488
rect 44177 39451 44235 39457
rect 45557 39457 45569 39460
rect 45603 39457 45615 39491
rect 45557 39451 45615 39457
rect 46477 39491 46535 39497
rect 46477 39457 46489 39491
rect 46523 39457 46535 39491
rect 46477 39451 46535 39457
rect 42852 39423 42883 39429
rect 42871 39389 42883 39423
rect 42852 39383 42883 39389
rect 43073 39423 43131 39429
rect 43073 39389 43085 39423
rect 43119 39389 43131 39423
rect 43073 39383 43131 39389
rect 42852 39380 42858 39383
rect 43162 39380 43168 39432
rect 43220 39429 43226 39432
rect 43220 39420 43228 39429
rect 44266 39420 44272 39432
rect 43220 39392 43265 39420
rect 44179 39392 44272 39420
rect 43220 39383 43228 39392
rect 43220 39380 43226 39383
rect 44266 39380 44272 39392
rect 44324 39420 44330 39432
rect 45649 39423 45707 39429
rect 44324 39392 45600 39420
rect 44324 39380 44330 39392
rect 45572 39364 45600 39392
rect 45649 39389 45661 39423
rect 45695 39389 45707 39423
rect 46934 39420 46940 39432
rect 46895 39392 46940 39420
rect 45649 39383 45707 39389
rect 41874 39352 41880 39364
rect 41386 39324 41644 39352
rect 41835 39324 41880 39352
rect 41141 39315 41199 39321
rect 34480 39256 36032 39284
rect 36817 39287 36875 39293
rect 34480 39244 34486 39256
rect 36817 39253 36829 39287
rect 36863 39284 36875 39287
rect 36906 39284 36912 39296
rect 36863 39256 36912 39284
rect 36863 39253 36875 39256
rect 36817 39247 36875 39253
rect 36906 39244 36912 39256
rect 36964 39244 36970 39296
rect 41156 39284 41184 39315
rect 41414 39284 41420 39296
rect 41156 39256 41420 39284
rect 41414 39244 41420 39256
rect 41472 39244 41478 39296
rect 41616 39293 41644 39324
rect 41874 39312 41880 39324
rect 41932 39312 41938 39364
rect 42978 39352 42984 39364
rect 42939 39324 42984 39352
rect 42978 39312 42984 39324
rect 43036 39312 43042 39364
rect 45554 39312 45560 39364
rect 45612 39312 45618 39364
rect 41601 39287 41659 39293
rect 41601 39253 41613 39287
rect 41647 39253 41659 39287
rect 41601 39247 41659 39253
rect 42426 39244 42432 39296
rect 42484 39284 42490 39296
rect 45462 39284 45468 39296
rect 42484 39256 45468 39284
rect 42484 39244 42490 39256
rect 45462 39244 45468 39256
rect 45520 39284 45526 39296
rect 45664 39284 45692 39383
rect 46934 39380 46940 39392
rect 46992 39380 46998 39432
rect 47026 39380 47032 39432
rect 47084 39420 47090 39432
rect 47228 39420 47256 39519
rect 49786 39516 49792 39528
rect 49844 39516 49850 39568
rect 52086 39516 52092 39568
rect 52144 39556 52150 39568
rect 53469 39559 53527 39565
rect 52144 39528 52960 39556
rect 52144 39516 52150 39528
rect 49694 39488 49700 39500
rect 48424 39460 49700 39488
rect 48041 39423 48099 39429
rect 48041 39420 48053 39423
rect 47084 39392 47129 39420
rect 47228 39392 48053 39420
rect 47084 39380 47090 39392
rect 48041 39389 48053 39392
rect 48087 39389 48099 39423
rect 48041 39383 48099 39389
rect 48189 39423 48247 39429
rect 48189 39389 48201 39423
rect 48235 39420 48247 39423
rect 48424 39420 48452 39460
rect 49694 39448 49700 39460
rect 49752 39488 49758 39500
rect 50341 39491 50399 39497
rect 50341 39488 50353 39491
rect 49752 39460 50353 39488
rect 49752 39448 49758 39460
rect 50341 39457 50353 39460
rect 50387 39457 50399 39491
rect 50341 39451 50399 39457
rect 51718 39448 51724 39500
rect 51776 39488 51782 39500
rect 52549 39491 52607 39497
rect 52549 39488 52561 39491
rect 51776 39460 52561 39488
rect 51776 39448 51782 39460
rect 52549 39457 52561 39460
rect 52595 39457 52607 39491
rect 52549 39451 52607 39457
rect 48235 39392 48452 39420
rect 48235 39389 48247 39392
rect 48189 39383 48247 39389
rect 48498 39380 48504 39432
rect 48556 39429 48562 39432
rect 48556 39420 48564 39429
rect 48866 39420 48872 39432
rect 48556 39392 48872 39420
rect 48556 39383 48564 39392
rect 48556 39380 48562 39383
rect 48866 39380 48872 39392
rect 48924 39380 48930 39432
rect 51092 39392 51764 39420
rect 47210 39352 47216 39364
rect 47171 39324 47216 39352
rect 47210 39312 47216 39324
rect 47268 39312 47274 39364
rect 48314 39352 48320 39364
rect 48275 39324 48320 39352
rect 48314 39312 48320 39324
rect 48372 39312 48378 39364
rect 48406 39312 48412 39364
rect 48464 39352 48470 39364
rect 49697 39355 49755 39361
rect 49697 39352 49709 39355
rect 48464 39324 48509 39352
rect 48613 39324 49709 39352
rect 48464 39312 48470 39324
rect 45520 39256 45692 39284
rect 45520 39244 45526 39256
rect 48130 39244 48136 39296
rect 48188 39284 48194 39296
rect 48613 39284 48641 39324
rect 49697 39321 49709 39324
rect 49743 39352 49755 39355
rect 50982 39352 50988 39364
rect 49743 39324 50988 39352
rect 49743 39321 49755 39324
rect 49697 39315 49755 39321
rect 50982 39312 50988 39324
rect 51040 39312 51046 39364
rect 48188 39256 48641 39284
rect 48188 39244 48194 39256
rect 48682 39244 48688 39296
rect 48740 39284 48746 39296
rect 49145 39287 49203 39293
rect 49145 39284 49157 39287
rect 48740 39256 49157 39284
rect 48740 39244 48746 39256
rect 49145 39253 49157 39256
rect 49191 39253 49203 39287
rect 49145 39247 49203 39253
rect 49326 39244 49332 39296
rect 49384 39284 49390 39296
rect 51092 39293 51120 39392
rect 51626 39352 51632 39364
rect 51587 39324 51632 39352
rect 51626 39312 51632 39324
rect 51684 39312 51690 39364
rect 51736 39352 51764 39392
rect 51810 39380 51816 39432
rect 51868 39420 51874 39432
rect 51905 39423 51963 39429
rect 51905 39420 51917 39423
rect 51868 39392 51917 39420
rect 51868 39380 51874 39392
rect 51905 39389 51917 39392
rect 51951 39389 51963 39423
rect 51905 39383 51963 39389
rect 51736 39324 51856 39352
rect 51077 39287 51135 39293
rect 51077 39284 51089 39287
rect 49384 39256 51089 39284
rect 49384 39244 49390 39256
rect 51077 39253 51089 39256
rect 51123 39253 51135 39287
rect 51718 39284 51724 39296
rect 51776 39293 51782 39296
rect 51828 39293 51856 39324
rect 51685 39256 51724 39284
rect 51077 39247 51135 39253
rect 51718 39244 51724 39256
rect 51776 39247 51785 39293
rect 51813 39287 51871 39293
rect 51813 39253 51825 39287
rect 51859 39284 51871 39287
rect 51902 39284 51908 39296
rect 51859 39256 51908 39284
rect 51859 39253 51871 39256
rect 51813 39247 51871 39253
rect 51776 39244 51782 39247
rect 51902 39244 51908 39256
rect 51960 39244 51966 39296
rect 52564 39284 52592 39451
rect 52932 39420 52960 39528
rect 53469 39525 53481 39559
rect 53515 39525 53527 39559
rect 53469 39519 53527 39525
rect 53374 39488 53380 39500
rect 53335 39460 53380 39488
rect 53374 39448 53380 39460
rect 53432 39448 53438 39500
rect 53285 39423 53343 39429
rect 53285 39420 53297 39423
rect 52932 39392 53297 39420
rect 53285 39389 53297 39392
rect 53331 39389 53343 39423
rect 53483 39420 53511 39519
rect 53561 39491 53619 39497
rect 53561 39457 53573 39491
rect 53607 39488 53619 39491
rect 53742 39488 53748 39500
rect 53607 39460 53748 39488
rect 53607 39457 53619 39460
rect 53561 39451 53619 39457
rect 53742 39448 53748 39460
rect 53800 39448 53806 39500
rect 53852 39488 53880 39596
rect 55677 39491 55735 39497
rect 55677 39488 55689 39491
rect 53852 39460 55689 39488
rect 55677 39457 55689 39460
rect 55723 39488 55735 39491
rect 55950 39488 55956 39500
rect 55723 39460 55956 39488
rect 55723 39457 55735 39460
rect 55677 39451 55735 39457
rect 55950 39448 55956 39460
rect 56008 39448 56014 39500
rect 54021 39423 54079 39429
rect 54021 39420 54033 39423
rect 53483 39392 54033 39420
rect 53285 39383 53343 39389
rect 54021 39389 54033 39392
rect 54067 39389 54079 39423
rect 54021 39383 54079 39389
rect 53300 39352 53328 39383
rect 54110 39380 54116 39432
rect 54168 39420 54174 39432
rect 54168 39392 54213 39420
rect 54168 39380 54174 39392
rect 54294 39380 54300 39432
rect 54352 39420 54358 39432
rect 54527 39423 54585 39429
rect 54352 39392 54397 39420
rect 54352 39380 54358 39392
rect 54527 39389 54539 39423
rect 54573 39420 54585 39423
rect 54754 39420 54760 39432
rect 54573 39392 54760 39420
rect 54573 39389 54585 39392
rect 54527 39383 54585 39389
rect 54754 39380 54760 39392
rect 54812 39380 54818 39432
rect 55766 39420 55772 39432
rect 55727 39392 55772 39420
rect 55766 39380 55772 39392
rect 55824 39380 55830 39432
rect 56870 39380 56876 39432
rect 56928 39420 56934 39432
rect 57057 39423 57115 39429
rect 57057 39420 57069 39423
rect 56928 39392 57069 39420
rect 56928 39380 56934 39392
rect 57057 39389 57069 39392
rect 57103 39389 57115 39423
rect 57238 39420 57244 39432
rect 57199 39392 57244 39420
rect 57057 39383 57115 39389
rect 57238 39380 57244 39392
rect 57296 39380 57302 39432
rect 54389 39355 54447 39361
rect 54389 39352 54401 39355
rect 53300 39324 54401 39352
rect 54128 39296 54156 39324
rect 54389 39321 54401 39324
rect 54435 39352 54447 39355
rect 55582 39352 55588 39364
rect 54435 39324 55588 39352
rect 54435 39321 54447 39324
rect 54389 39315 54447 39321
rect 55582 39312 55588 39324
rect 55640 39312 55646 39364
rect 53466 39284 53472 39296
rect 52564 39256 53472 39284
rect 53466 39244 53472 39256
rect 53524 39244 53530 39296
rect 54110 39244 54116 39296
rect 54168 39244 54174 39296
rect 54665 39287 54723 39293
rect 54665 39253 54677 39287
rect 54711 39284 54723 39287
rect 56042 39284 56048 39296
rect 54711 39256 56048 39284
rect 54711 39253 54723 39256
rect 54665 39247 54723 39253
rect 56042 39244 56048 39256
rect 56100 39244 56106 39296
rect 56137 39287 56195 39293
rect 56137 39253 56149 39287
rect 56183 39284 56195 39287
rect 56502 39284 56508 39296
rect 56183 39256 56508 39284
rect 56183 39253 56195 39256
rect 56137 39247 56195 39253
rect 56502 39244 56508 39256
rect 56560 39244 56566 39296
rect 58069 39287 58127 39293
rect 58069 39253 58081 39287
rect 58115 39284 58127 39287
rect 58434 39284 58440 39296
rect 58115 39256 58440 39284
rect 58115 39253 58127 39256
rect 58069 39247 58127 39253
rect 58434 39244 58440 39256
rect 58492 39244 58498 39296
rect 1104 39194 58880 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 35594 39194
rect 35646 39142 35658 39194
rect 35710 39142 35722 39194
rect 35774 39142 35786 39194
rect 35838 39142 35850 39194
rect 35902 39142 58880 39194
rect 1104 39120 58880 39142
rect 30558 39080 30564 39092
rect 30519 39052 30564 39080
rect 30558 39040 30564 39052
rect 30616 39040 30622 39092
rect 31573 39083 31631 39089
rect 31573 39049 31585 39083
rect 31619 39080 31631 39083
rect 31662 39080 31668 39092
rect 31619 39052 31668 39080
rect 31619 39049 31631 39052
rect 31573 39043 31631 39049
rect 31662 39040 31668 39052
rect 31720 39040 31726 39092
rect 32490 39040 32496 39092
rect 32548 39080 32554 39092
rect 32861 39083 32919 39089
rect 32861 39080 32873 39083
rect 32548 39052 32873 39080
rect 32548 39040 32554 39052
rect 32861 39049 32873 39052
rect 32907 39049 32919 39083
rect 34422 39080 34428 39092
rect 34383 39052 34428 39080
rect 32861 39043 32919 39049
rect 32766 39012 32772 39024
rect 31496 38984 32772 39012
rect 29730 38944 29736 38956
rect 29691 38916 29736 38944
rect 29730 38904 29736 38916
rect 29788 38904 29794 38956
rect 30745 38947 30803 38953
rect 30745 38913 30757 38947
rect 30791 38944 30803 38947
rect 30834 38944 30840 38956
rect 30791 38916 30840 38944
rect 30791 38913 30803 38916
rect 30745 38907 30803 38913
rect 30834 38904 30840 38916
rect 30892 38904 30898 38956
rect 31496 38953 31524 38984
rect 32766 38972 32772 38984
rect 32824 38972 32830 39024
rect 32876 39012 32904 39043
rect 34422 39040 34428 39052
rect 34480 39040 34486 39092
rect 35434 39040 35440 39092
rect 35492 39080 35498 39092
rect 35529 39083 35587 39089
rect 35529 39080 35541 39083
rect 35492 39052 35541 39080
rect 35492 39040 35498 39052
rect 35529 39049 35541 39052
rect 35575 39049 35587 39083
rect 35529 39043 35587 39049
rect 41969 39083 42027 39089
rect 41969 39049 41981 39083
rect 42015 39080 42027 39083
rect 44266 39080 44272 39092
rect 42015 39052 44272 39080
rect 42015 39049 42027 39052
rect 41969 39043 42027 39049
rect 44266 39040 44272 39052
rect 44324 39040 44330 39092
rect 46293 39083 46351 39089
rect 46293 39049 46305 39083
rect 46339 39080 46351 39083
rect 47026 39080 47032 39092
rect 46339 39052 47032 39080
rect 46339 39049 46351 39052
rect 46293 39043 46351 39049
rect 47026 39040 47032 39052
rect 47084 39040 47090 39092
rect 47121 39083 47179 39089
rect 47121 39049 47133 39083
rect 47167 39080 47179 39083
rect 47578 39080 47584 39092
rect 47167 39052 47584 39080
rect 47167 39049 47179 39052
rect 47121 39043 47179 39049
rect 47578 39040 47584 39052
rect 47636 39040 47642 39092
rect 48406 39080 48412 39092
rect 48056 39052 48412 39080
rect 36538 39012 36544 39024
rect 32876 38984 35388 39012
rect 36499 38984 36544 39012
rect 31481 38947 31539 38953
rect 31481 38913 31493 38947
rect 31527 38913 31539 38947
rect 31757 38947 31815 38953
rect 31757 38944 31769 38947
rect 31481 38907 31539 38913
rect 31588 38916 31769 38944
rect 29178 38836 29184 38888
rect 29236 38876 29242 38888
rect 30009 38879 30067 38885
rect 30009 38876 30021 38879
rect 29236 38848 30021 38876
rect 29236 38836 29242 38848
rect 30009 38845 30021 38848
rect 30055 38876 30067 38879
rect 31496 38876 31524 38907
rect 30055 38848 31524 38876
rect 30055 38845 30067 38848
rect 30009 38839 30067 38845
rect 29825 38811 29883 38817
rect 29825 38777 29837 38811
rect 29871 38808 29883 38811
rect 31588 38808 31616 38916
rect 31757 38913 31769 38916
rect 31803 38944 31815 38947
rect 32306 38944 32312 38956
rect 31803 38916 32312 38944
rect 31803 38913 31815 38916
rect 31757 38907 31815 38913
rect 32306 38904 32312 38916
rect 32364 38904 32370 38956
rect 32674 38904 32680 38956
rect 32732 38944 32738 38956
rect 32953 38947 33011 38953
rect 32953 38944 32965 38947
rect 32732 38916 32965 38944
rect 32732 38904 32738 38916
rect 32953 38913 32965 38916
rect 32999 38913 33011 38947
rect 32953 38907 33011 38913
rect 33594 38904 33600 38956
rect 33652 38944 33658 38956
rect 34057 38947 34115 38953
rect 34057 38944 34069 38947
rect 33652 38916 34069 38944
rect 33652 38904 33658 38916
rect 34057 38913 34069 38916
rect 34103 38913 34115 38947
rect 34057 38907 34115 38913
rect 34606 38904 34612 38956
rect 34664 38944 34670 38956
rect 35250 38944 35256 38956
rect 34664 38916 35256 38944
rect 34664 38904 34670 38916
rect 35250 38904 35256 38916
rect 35308 38904 35314 38956
rect 35360 38944 35388 38984
rect 36538 38972 36544 38984
rect 36596 38972 36602 39024
rect 41414 38972 41420 39024
rect 41472 39012 41478 39024
rect 42426 39012 42432 39024
rect 41472 38984 42432 39012
rect 41472 38972 41478 38984
rect 42426 38972 42432 38984
rect 42484 38972 42490 39024
rect 45097 39015 45155 39021
rect 45097 39012 45109 39015
rect 42628 38984 45109 39012
rect 36403 38947 36461 38953
rect 36403 38944 36415 38947
rect 35360 38916 36415 38944
rect 36403 38913 36415 38916
rect 36449 38913 36461 38947
rect 36633 38947 36691 38953
rect 36633 38944 36645 38947
rect 36403 38907 36461 38913
rect 36556 38916 36645 38944
rect 33870 38836 33876 38888
rect 33928 38876 33934 38888
rect 33965 38879 34023 38885
rect 33965 38876 33977 38879
rect 33928 38848 33977 38876
rect 33928 38836 33934 38848
rect 33965 38845 33977 38848
rect 34011 38845 34023 38879
rect 33965 38839 34023 38845
rect 34698 38836 34704 38888
rect 34756 38876 34762 38888
rect 35342 38876 35348 38888
rect 34756 38848 35348 38876
rect 34756 38836 34762 38848
rect 35342 38836 35348 38848
rect 35400 38836 35406 38888
rect 35434 38836 35440 38888
rect 35492 38876 35498 38888
rect 35529 38879 35587 38885
rect 35529 38876 35541 38879
rect 35492 38848 35541 38876
rect 35492 38836 35498 38848
rect 35529 38845 35541 38848
rect 35575 38845 35587 38879
rect 35529 38839 35587 38845
rect 29871 38780 31616 38808
rect 29871 38777 29883 38780
rect 29825 38771 29883 38777
rect 33042 38768 33048 38820
rect 33100 38808 33106 38820
rect 36556 38808 36584 38916
rect 36633 38913 36645 38916
rect 36679 38913 36691 38947
rect 36814 38944 36820 38956
rect 36775 38916 36820 38944
rect 36633 38907 36691 38913
rect 36814 38904 36820 38916
rect 36872 38904 36878 38956
rect 36906 38904 36912 38956
rect 36964 38944 36970 38956
rect 36964 38916 37009 38944
rect 36964 38904 36970 38916
rect 38102 38904 38108 38956
rect 38160 38944 38166 38956
rect 38565 38947 38623 38953
rect 38565 38944 38577 38947
rect 38160 38916 38577 38944
rect 38160 38904 38166 38916
rect 38565 38913 38577 38916
rect 38611 38913 38623 38947
rect 38565 38907 38623 38913
rect 38654 38904 38660 38956
rect 38712 38944 38718 38956
rect 39209 38947 39267 38953
rect 39209 38944 39221 38947
rect 38712 38916 39221 38944
rect 38712 38904 38718 38916
rect 39209 38913 39221 38916
rect 39255 38913 39267 38947
rect 39209 38907 39267 38913
rect 40034 38904 40040 38956
rect 40092 38944 40098 38956
rect 42628 38953 42656 38984
rect 45097 38981 45109 38984
rect 45143 38981 45155 39015
rect 45097 38975 45155 38981
rect 41141 38947 41199 38953
rect 41141 38944 41153 38947
rect 40092 38916 41153 38944
rect 40092 38904 40098 38916
rect 41141 38913 41153 38916
rect 41187 38913 41199 38947
rect 41141 38907 41199 38913
rect 42613 38947 42671 38953
rect 42613 38913 42625 38947
rect 42659 38913 42671 38947
rect 42613 38907 42671 38913
rect 42706 38947 42764 38953
rect 42706 38913 42718 38947
rect 42752 38913 42764 38947
rect 42886 38944 42892 38956
rect 42847 38916 42892 38944
rect 42706 38907 42764 38913
rect 39850 38876 39856 38888
rect 39811 38848 39856 38876
rect 39850 38836 39856 38848
rect 39908 38836 39914 38888
rect 41046 38876 41052 38888
rect 41007 38848 41052 38876
rect 41046 38836 41052 38848
rect 41104 38836 41110 38888
rect 37734 38808 37740 38820
rect 33100 38780 37740 38808
rect 33100 38768 33106 38780
rect 37734 38768 37740 38780
rect 37792 38768 37798 38820
rect 41156 38808 41184 38907
rect 41966 38836 41972 38888
rect 42024 38876 42030 38888
rect 42720 38876 42748 38907
rect 42886 38904 42892 38916
rect 42944 38904 42950 38956
rect 43162 38953 43168 38956
rect 42981 38947 43039 38953
rect 42981 38913 42993 38947
rect 43027 38913 43039 38947
rect 42981 38907 43039 38913
rect 43119 38947 43168 38953
rect 43119 38913 43131 38947
rect 43165 38913 43168 38947
rect 43119 38907 43168 38913
rect 42024 38848 42748 38876
rect 42024 38836 42030 38848
rect 42794 38836 42800 38888
rect 42852 38876 42858 38888
rect 42996 38876 43024 38907
rect 43162 38904 43168 38907
rect 43220 38904 43226 38956
rect 44174 38944 44180 38956
rect 44135 38916 44180 38944
rect 44174 38904 44180 38916
rect 44232 38904 44238 38956
rect 45002 38944 45008 38956
rect 44963 38916 45008 38944
rect 45002 38904 45008 38916
rect 45060 38904 45066 38956
rect 45186 38944 45192 38956
rect 45147 38916 45192 38944
rect 45186 38904 45192 38916
rect 45244 38904 45250 38956
rect 46477 38947 46535 38953
rect 46477 38913 46489 38947
rect 46523 38913 46535 38947
rect 46477 38907 46535 38913
rect 46937 38947 46995 38953
rect 46937 38913 46949 38947
rect 46983 38944 46995 38947
rect 48056 38944 48084 39052
rect 48406 39040 48412 39052
rect 48464 39080 48470 39092
rect 48866 39080 48872 39092
rect 48464 39052 48636 39080
rect 48464 39040 48470 39052
rect 48130 38972 48136 39024
rect 48188 39012 48194 39024
rect 48608 39021 48636 39052
rect 48792 39052 48872 39080
rect 48593 39015 48651 39021
rect 48188 38984 48453 39012
rect 48188 38972 48194 38984
rect 48314 38944 48320 38956
rect 46983 38916 48084 38944
rect 48275 38916 48320 38944
rect 46983 38913 46995 38916
rect 46937 38907 46995 38913
rect 44085 38879 44143 38885
rect 44085 38876 44097 38879
rect 42852 38848 43024 38876
rect 43272 38848 44097 38876
rect 42852 38836 42858 38848
rect 43272 38817 43300 38848
rect 44085 38845 44097 38848
rect 44131 38845 44143 38879
rect 46492 38876 46520 38907
rect 48314 38904 48320 38916
rect 48372 38904 48378 38956
rect 48425 38953 48453 38984
rect 48593 38981 48605 39015
rect 48639 38981 48651 39015
rect 48593 38975 48651 38981
rect 48792 38953 48820 39052
rect 48866 39040 48872 39052
rect 48924 39040 48930 39092
rect 48961 39083 49019 39089
rect 48961 39049 48973 39083
rect 49007 39080 49019 39083
rect 55766 39080 55772 39092
rect 49007 39052 55772 39080
rect 49007 39049 49019 39052
rect 48961 39043 49019 39049
rect 55766 39040 55772 39052
rect 55824 39040 55830 39092
rect 56870 39080 56876 39092
rect 56831 39052 56876 39080
rect 56870 39040 56876 39052
rect 56928 39040 56934 39092
rect 50249 39015 50307 39021
rect 50249 39012 50261 39015
rect 48884 38984 50261 39012
rect 48410 38947 48468 38953
rect 48410 38913 48422 38947
rect 48456 38913 48468 38947
rect 48410 38907 48468 38913
rect 48685 38947 48743 38953
rect 48685 38913 48697 38947
rect 48731 38913 48743 38947
rect 48685 38907 48743 38913
rect 48782 38947 48840 38953
rect 48782 38913 48794 38947
rect 48828 38913 48840 38947
rect 48782 38907 48840 38913
rect 47210 38876 47216 38888
rect 46492 38848 47216 38876
rect 44085 38839 44143 38845
rect 47210 38836 47216 38848
rect 47268 38876 47274 38888
rect 47762 38876 47768 38888
rect 47268 38848 47768 38876
rect 47268 38836 47274 38848
rect 47762 38836 47768 38848
rect 47820 38836 47826 38888
rect 47854 38836 47860 38888
rect 47912 38876 47918 38888
rect 47912 38848 48452 38876
rect 47912 38836 47918 38848
rect 43257 38811 43315 38817
rect 41156 38780 42840 38808
rect 29917 38743 29975 38749
rect 29917 38709 29929 38743
rect 29963 38740 29975 38743
rect 30374 38740 30380 38752
rect 29963 38712 30380 38740
rect 29963 38709 29975 38712
rect 29917 38703 29975 38709
rect 30374 38700 30380 38712
rect 30432 38700 30438 38752
rect 31757 38743 31815 38749
rect 31757 38709 31769 38743
rect 31803 38740 31815 38743
rect 32214 38740 32220 38752
rect 31803 38712 32220 38740
rect 31803 38709 31815 38712
rect 31757 38703 31815 38709
rect 32214 38700 32220 38712
rect 32272 38700 32278 38752
rect 36265 38743 36323 38749
rect 36265 38709 36277 38743
rect 36311 38740 36323 38743
rect 37274 38740 37280 38752
rect 36311 38712 37280 38740
rect 36311 38709 36323 38712
rect 36265 38703 36323 38709
rect 37274 38700 37280 38712
rect 37332 38700 37338 38752
rect 37550 38740 37556 38752
rect 37511 38712 37556 38740
rect 37550 38700 37556 38712
rect 37608 38700 37614 38752
rect 42058 38700 42064 38752
rect 42116 38740 42122 38752
rect 42702 38740 42708 38752
rect 42116 38712 42708 38740
rect 42116 38700 42122 38712
rect 42702 38700 42708 38712
rect 42760 38700 42766 38752
rect 42812 38740 42840 38780
rect 43257 38777 43269 38811
rect 43303 38777 43315 38811
rect 43257 38771 43315 38777
rect 44545 38811 44603 38817
rect 44545 38777 44557 38811
rect 44591 38808 44603 38811
rect 45738 38808 45744 38820
rect 44591 38780 45744 38808
rect 44591 38777 44603 38780
rect 44545 38771 44603 38777
rect 45738 38768 45744 38780
rect 45796 38768 45802 38820
rect 47118 38768 47124 38820
rect 47176 38808 47182 38820
rect 48424 38808 48452 38848
rect 48700 38808 48728 38907
rect 47176 38780 48360 38808
rect 48424 38780 48728 38808
rect 47176 38768 47182 38780
rect 43806 38740 43812 38752
rect 42812 38712 43812 38740
rect 43806 38700 43812 38712
rect 43864 38700 43870 38752
rect 45646 38740 45652 38752
rect 45607 38712 45652 38740
rect 45646 38700 45652 38712
rect 45704 38700 45710 38752
rect 47854 38740 47860 38752
rect 47815 38712 47860 38740
rect 47854 38700 47860 38712
rect 47912 38700 47918 38752
rect 48332 38740 48360 38780
rect 48884 38740 48912 38984
rect 50249 38981 50261 38984
rect 50295 39012 50307 39015
rect 51626 39012 51632 39024
rect 50295 38984 51632 39012
rect 50295 38981 50307 38984
rect 50249 38975 50307 38981
rect 51626 38972 51632 38984
rect 51684 38972 51690 39024
rect 51718 38972 51724 39024
rect 51776 39012 51782 39024
rect 51776 38984 53604 39012
rect 51776 38972 51782 38984
rect 49050 38904 49056 38956
rect 49108 38944 49114 38956
rect 49973 38947 50031 38953
rect 49973 38944 49985 38947
rect 49108 38916 49985 38944
rect 49108 38904 49114 38916
rect 49973 38913 49985 38916
rect 50019 38913 50031 38947
rect 49973 38907 50031 38913
rect 50065 38947 50123 38953
rect 50065 38913 50077 38947
rect 50111 38944 50123 38947
rect 50706 38944 50712 38956
rect 50111 38916 50712 38944
rect 50111 38913 50123 38916
rect 50065 38907 50123 38913
rect 49988 38808 50016 38907
rect 50706 38904 50712 38916
rect 50764 38904 50770 38956
rect 51074 38904 51080 38956
rect 51132 38944 51138 38956
rect 51132 38916 51177 38944
rect 51132 38904 51138 38916
rect 51994 38904 52000 38956
rect 52052 38904 52058 38956
rect 52822 38904 52828 38956
rect 52880 38944 52886 38956
rect 53055 38947 53113 38953
rect 53055 38944 53067 38947
rect 52880 38916 53067 38944
rect 52880 38904 52886 38916
rect 53055 38913 53067 38916
rect 53101 38913 53113 38947
rect 53055 38907 53113 38913
rect 53193 38947 53251 38953
rect 53193 38913 53205 38947
rect 53239 38913 53251 38947
rect 53193 38907 53251 38913
rect 53285 38947 53343 38953
rect 53285 38913 53297 38947
rect 53331 38913 53343 38947
rect 53466 38944 53472 38956
rect 53427 38916 53472 38944
rect 53285 38907 53343 38913
rect 51166 38876 51172 38888
rect 51127 38848 51172 38876
rect 51166 38836 51172 38848
rect 51224 38836 51230 38888
rect 51905 38879 51963 38885
rect 51905 38845 51917 38879
rect 51951 38845 51963 38879
rect 52012 38876 52040 38904
rect 53208 38876 53236 38907
rect 52012 38848 53236 38876
rect 51905 38839 51963 38845
rect 50798 38808 50804 38820
rect 49988 38780 50804 38808
rect 50798 38768 50804 38780
rect 50856 38808 50862 38820
rect 51810 38808 51816 38820
rect 50856 38780 51816 38808
rect 50856 38768 50862 38780
rect 51810 38768 51816 38780
rect 51868 38768 51874 38820
rect 48332 38712 48912 38740
rect 49326 38700 49332 38752
rect 49384 38740 49390 38752
rect 49421 38743 49479 38749
rect 49421 38740 49433 38743
rect 49384 38712 49433 38740
rect 49384 38700 49390 38712
rect 49421 38709 49433 38712
rect 49467 38709 49479 38743
rect 49421 38703 49479 38709
rect 50249 38743 50307 38749
rect 50249 38709 50261 38743
rect 50295 38740 50307 38743
rect 50338 38740 50344 38752
rect 50295 38712 50344 38740
rect 50295 38709 50307 38712
rect 50249 38703 50307 38709
rect 50338 38700 50344 38712
rect 50396 38700 50402 38752
rect 51920 38740 51948 38839
rect 51994 38768 52000 38820
rect 52052 38808 52058 38820
rect 52270 38808 52276 38820
rect 52052 38780 52276 38808
rect 52052 38768 52058 38780
rect 52270 38768 52276 38780
rect 52328 38808 52334 38820
rect 53300 38808 53328 38907
rect 53466 38904 53472 38916
rect 53524 38904 53530 38956
rect 53576 38953 53604 38984
rect 54110 38972 54116 39024
rect 54168 39012 54174 39024
rect 54168 38984 54341 39012
rect 54168 38972 54174 38984
rect 53561 38947 53619 38953
rect 53561 38913 53573 38947
rect 53607 38913 53619 38947
rect 54202 38944 54208 38956
rect 54163 38916 54208 38944
rect 53561 38907 53619 38913
rect 54202 38904 54208 38916
rect 54260 38904 54266 38956
rect 54313 38953 54341 38984
rect 54386 38972 54392 39024
rect 54444 39012 54450 39024
rect 54481 39015 54539 39021
rect 54481 39012 54493 39015
rect 54444 38984 54493 39012
rect 54444 38972 54450 38984
rect 54481 38981 54493 38984
rect 54527 38981 54539 39015
rect 54481 38975 54539 38981
rect 54298 38947 54356 38953
rect 54298 38913 54310 38947
rect 54344 38913 54356 38947
rect 54298 38907 54356 38913
rect 54573 38947 54631 38953
rect 54573 38913 54585 38947
rect 54619 38913 54631 38947
rect 54573 38907 54631 38913
rect 53484 38876 53512 38904
rect 53834 38876 53840 38888
rect 53484 38848 53840 38876
rect 53834 38836 53840 38848
rect 53892 38836 53898 38888
rect 54018 38836 54024 38888
rect 54076 38876 54082 38888
rect 54588 38876 54616 38907
rect 54662 38904 54668 38956
rect 54720 38953 54726 38956
rect 54720 38944 54728 38953
rect 56502 38944 56508 38956
rect 54720 38916 54765 38944
rect 56463 38916 56508 38944
rect 54720 38907 54728 38916
rect 54720 38904 54726 38907
rect 56502 38904 56508 38916
rect 56560 38904 56566 38956
rect 55309 38879 55367 38885
rect 55309 38876 55321 38879
rect 54076 38848 55321 38876
rect 54076 38836 54082 38848
rect 55309 38845 55321 38848
rect 55355 38845 55367 38879
rect 55309 38839 55367 38845
rect 52328 38780 53328 38808
rect 55324 38808 55352 38839
rect 56042 38836 56048 38888
rect 56100 38876 56106 38888
rect 56413 38879 56471 38885
rect 56413 38876 56425 38879
rect 56100 38848 56425 38876
rect 56100 38836 56106 38848
rect 56413 38845 56425 38848
rect 56459 38845 56471 38879
rect 56413 38839 56471 38845
rect 57333 38811 57391 38817
rect 57333 38808 57345 38811
rect 55324 38780 57345 38808
rect 52328 38768 52334 38780
rect 57333 38777 57345 38780
rect 57379 38777 57391 38811
rect 57333 38771 57391 38777
rect 52730 38740 52736 38752
rect 51920 38712 52736 38740
rect 52730 38700 52736 38712
rect 52788 38700 52794 38752
rect 52917 38743 52975 38749
rect 52917 38709 52929 38743
rect 52963 38740 52975 38743
rect 53006 38740 53012 38752
rect 52963 38712 53012 38740
rect 52963 38709 52975 38712
rect 52917 38703 52975 38709
rect 53006 38700 53012 38712
rect 53064 38700 53070 38752
rect 54849 38743 54907 38749
rect 54849 38709 54861 38743
rect 54895 38740 54907 38743
rect 55214 38740 55220 38752
rect 54895 38712 55220 38740
rect 54895 38709 54907 38712
rect 54849 38703 54907 38709
rect 55214 38700 55220 38712
rect 55272 38700 55278 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 30650 38496 30656 38548
rect 30708 38536 30714 38548
rect 31297 38539 31355 38545
rect 31297 38536 31309 38539
rect 30708 38508 31309 38536
rect 30708 38496 30714 38508
rect 31297 38505 31309 38508
rect 31343 38505 31355 38539
rect 33870 38536 33876 38548
rect 31297 38499 31355 38505
rect 31726 38508 32996 38536
rect 33831 38508 33876 38536
rect 28997 38471 29055 38477
rect 28997 38437 29009 38471
rect 29043 38437 29055 38471
rect 31726 38468 31754 38508
rect 28997 38431 29055 38437
rect 31036 38440 31754 38468
rect 29012 38400 29040 38431
rect 31036 38400 31064 38440
rect 31846 38428 31852 38480
rect 31904 38468 31910 38480
rect 32861 38471 32919 38477
rect 31904 38440 32444 38468
rect 31904 38428 31910 38440
rect 29012 38372 31064 38400
rect 29181 38335 29239 38341
rect 29181 38301 29193 38335
rect 29227 38332 29239 38335
rect 30098 38332 30104 38344
rect 29227 38304 30104 38332
rect 29227 38301 29239 38304
rect 29181 38295 29239 38301
rect 30098 38292 30104 38304
rect 30156 38292 30162 38344
rect 30374 38292 30380 38344
rect 30432 38332 30438 38344
rect 31036 38341 31064 38372
rect 31202 38341 31208 38344
rect 30653 38335 30711 38341
rect 30653 38332 30665 38335
rect 30432 38304 30665 38332
rect 30432 38292 30438 38304
rect 30653 38301 30665 38304
rect 30699 38301 30711 38335
rect 30653 38295 30711 38301
rect 30801 38335 30859 38341
rect 30801 38301 30813 38335
rect 30847 38332 30859 38335
rect 31021 38335 31079 38341
rect 30847 38301 30880 38332
rect 30801 38295 30880 38301
rect 31021 38301 31033 38335
rect 31067 38301 31079 38335
rect 31021 38295 31079 38301
rect 31159 38335 31208 38341
rect 31159 38301 31171 38335
rect 31205 38301 31208 38335
rect 31159 38295 31208 38301
rect 29730 38224 29736 38276
rect 29788 38264 29794 38276
rect 29825 38267 29883 38273
rect 29825 38264 29837 38267
rect 29788 38236 29837 38264
rect 29788 38224 29794 38236
rect 29825 38233 29837 38236
rect 29871 38233 29883 38267
rect 29825 38227 29883 38233
rect 30101 38199 30159 38205
rect 30101 38165 30113 38199
rect 30147 38196 30159 38199
rect 30742 38196 30748 38208
rect 30147 38168 30748 38196
rect 30147 38165 30159 38168
rect 30101 38159 30159 38165
rect 30742 38156 30748 38168
rect 30800 38196 30806 38208
rect 30852 38196 30880 38295
rect 31202 38292 31208 38295
rect 31260 38292 31266 38344
rect 32214 38332 32220 38344
rect 32175 38304 32220 38332
rect 32214 38292 32220 38304
rect 32272 38292 32278 38344
rect 32310 38335 32368 38341
rect 32310 38301 32322 38335
rect 32356 38301 32368 38335
rect 32310 38295 32368 38301
rect 30929 38267 30987 38273
rect 30929 38233 30941 38267
rect 30975 38264 30987 38267
rect 31570 38264 31576 38276
rect 30975 38236 31576 38264
rect 30975 38233 30987 38236
rect 30929 38227 30987 38233
rect 31570 38224 31576 38236
rect 31628 38224 31634 38276
rect 31662 38224 31668 38276
rect 31720 38264 31726 38276
rect 32324 38264 32352 38295
rect 31720 38236 32352 38264
rect 32416 38264 32444 38440
rect 32861 38437 32873 38471
rect 32907 38437 32919 38471
rect 32968 38468 32996 38508
rect 33870 38496 33876 38508
rect 33928 38496 33934 38548
rect 35342 38536 35348 38548
rect 35303 38508 35348 38536
rect 35342 38496 35348 38508
rect 35400 38496 35406 38548
rect 35434 38496 35440 38548
rect 35492 38536 35498 38548
rect 35897 38539 35955 38545
rect 35897 38536 35909 38539
rect 35492 38508 35909 38536
rect 35492 38496 35498 38508
rect 35897 38505 35909 38508
rect 35943 38505 35955 38539
rect 41046 38536 41052 38548
rect 41007 38508 41052 38536
rect 35897 38499 35955 38505
rect 41046 38496 41052 38508
rect 41104 38496 41110 38548
rect 47210 38536 47216 38548
rect 47171 38508 47216 38536
rect 47210 38496 47216 38508
rect 47268 38496 47274 38548
rect 48133 38539 48191 38545
rect 48133 38505 48145 38539
rect 48179 38536 48191 38539
rect 48314 38536 48320 38548
rect 48179 38508 48320 38536
rect 48179 38505 48191 38508
rect 48133 38499 48191 38505
rect 48314 38496 48320 38508
rect 48372 38496 48378 38548
rect 50985 38539 51043 38545
rect 50985 38505 50997 38539
rect 51031 38536 51043 38539
rect 51074 38536 51080 38548
rect 51031 38508 51080 38536
rect 51031 38505 51043 38508
rect 50985 38499 51043 38505
rect 51074 38496 51080 38508
rect 51132 38496 51138 38548
rect 51902 38496 51908 38548
rect 51960 38536 51966 38548
rect 51997 38539 52055 38545
rect 51997 38536 52009 38539
rect 51960 38508 52009 38536
rect 51960 38496 51966 38508
rect 51997 38505 52009 38508
rect 52043 38505 52055 38539
rect 51997 38499 52055 38505
rect 52914 38496 52920 38548
rect 52972 38536 52978 38548
rect 53466 38536 53472 38548
rect 52972 38508 53472 38536
rect 52972 38496 52978 38508
rect 53466 38496 53472 38508
rect 53524 38536 53530 38548
rect 53929 38539 53987 38545
rect 53929 38536 53941 38539
rect 53524 38508 53941 38536
rect 53524 38496 53530 38508
rect 53929 38505 53941 38508
rect 53975 38505 53987 38539
rect 53929 38499 53987 38505
rect 54021 38539 54079 38545
rect 54021 38505 54033 38539
rect 54067 38536 54079 38539
rect 54202 38536 54208 38548
rect 54067 38508 54208 38536
rect 54067 38505 54079 38508
rect 54021 38499 54079 38505
rect 54202 38496 54208 38508
rect 54260 38496 54266 38548
rect 55306 38496 55312 38548
rect 55364 38536 55370 38548
rect 55582 38536 55588 38548
rect 55364 38508 55588 38536
rect 55364 38496 55370 38508
rect 55582 38496 55588 38508
rect 55640 38536 55646 38548
rect 56505 38539 56563 38545
rect 56505 38536 56517 38539
rect 55640 38508 56517 38536
rect 55640 38496 55646 38508
rect 56505 38505 56517 38508
rect 56551 38505 56563 38539
rect 56505 38499 56563 38505
rect 34606 38468 34612 38480
rect 32968 38440 34612 38468
rect 32861 38431 32919 38437
rect 32490 38292 32496 38344
rect 32548 38332 32554 38344
rect 32548 38304 32593 38332
rect 32548 38292 32554 38304
rect 32674 38292 32680 38344
rect 32732 38341 32738 38344
rect 32732 38332 32740 38341
rect 32876 38332 32904 38431
rect 34606 38428 34612 38440
rect 34664 38428 34670 38480
rect 36722 38468 36728 38480
rect 34808 38440 36728 38468
rect 33410 38400 33416 38412
rect 33371 38372 33416 38400
rect 33410 38360 33416 38372
rect 33468 38400 33474 38412
rect 33686 38400 33692 38412
rect 33468 38372 33692 38400
rect 33468 38360 33474 38372
rect 33686 38360 33692 38372
rect 33744 38360 33750 38412
rect 34808 38400 34836 38440
rect 36722 38428 36728 38440
rect 36780 38428 36786 38480
rect 40034 38468 40040 38480
rect 37936 38440 40040 38468
rect 36740 38400 36768 38428
rect 34440 38372 34836 38400
rect 34900 38372 36032 38400
rect 36740 38372 37780 38400
rect 33505 38335 33563 38341
rect 33505 38332 33517 38335
rect 32732 38304 32777 38332
rect 32876 38304 33517 38332
rect 32732 38295 32740 38304
rect 33505 38301 33517 38304
rect 33551 38301 33563 38335
rect 33505 38295 33563 38301
rect 32732 38292 32738 38295
rect 32585 38267 32643 38273
rect 32585 38264 32597 38267
rect 32416 38236 32597 38264
rect 31720 38224 31726 38236
rect 32585 38233 32597 38236
rect 32631 38264 32643 38267
rect 34440 38264 34468 38372
rect 34514 38292 34520 38344
rect 34572 38332 34578 38344
rect 34900 38341 34928 38372
rect 34885 38335 34943 38341
rect 34885 38332 34897 38335
rect 34572 38304 34897 38332
rect 34572 38292 34578 38304
rect 34885 38301 34897 38304
rect 34931 38301 34943 38335
rect 35066 38332 35072 38344
rect 35027 38304 35072 38332
rect 34885 38295 34943 38301
rect 35066 38292 35072 38304
rect 35124 38292 35130 38344
rect 36004 38341 36032 38372
rect 35897 38335 35955 38341
rect 35897 38301 35909 38335
rect 35943 38301 35955 38335
rect 35897 38295 35955 38301
rect 35989 38335 36047 38341
rect 35989 38301 36001 38335
rect 36035 38332 36047 38335
rect 36354 38332 36360 38344
rect 36035 38304 36360 38332
rect 36035 38301 36047 38304
rect 35989 38295 36047 38301
rect 32631 38236 34468 38264
rect 32631 38233 32643 38236
rect 32585 38227 32643 38233
rect 34974 38224 34980 38276
rect 35032 38264 35038 38276
rect 35437 38267 35495 38273
rect 35437 38264 35449 38267
rect 35032 38236 35449 38264
rect 35032 38224 35038 38236
rect 35437 38233 35449 38236
rect 35483 38264 35495 38267
rect 35912 38264 35940 38295
rect 36354 38292 36360 38304
rect 36412 38292 36418 38344
rect 36630 38332 36636 38344
rect 36464 38304 36636 38332
rect 35483 38236 35940 38264
rect 36173 38267 36231 38273
rect 35483 38233 35495 38236
rect 35437 38227 35495 38233
rect 36173 38233 36185 38267
rect 36219 38264 36231 38267
rect 36464 38264 36492 38304
rect 36630 38292 36636 38304
rect 36688 38292 36694 38344
rect 36814 38332 36820 38344
rect 36775 38304 36820 38332
rect 36814 38292 36820 38304
rect 36872 38292 36878 38344
rect 37274 38292 37280 38344
rect 37332 38332 37338 38344
rect 37553 38335 37611 38341
rect 37553 38332 37565 38335
rect 37332 38304 37565 38332
rect 37332 38292 37338 38304
rect 37553 38301 37565 38304
rect 37599 38301 37611 38335
rect 37553 38295 37611 38301
rect 36219 38236 36492 38264
rect 37752 38264 37780 38372
rect 37936 38344 37964 38440
rect 40034 38428 40040 38440
rect 40092 38428 40098 38480
rect 43901 38471 43959 38477
rect 43901 38437 43913 38471
rect 43947 38468 43959 38471
rect 44174 38468 44180 38480
rect 43947 38440 44180 38468
rect 43947 38437 43959 38440
rect 43901 38431 43959 38437
rect 44174 38428 44180 38440
rect 44232 38428 44238 38480
rect 49697 38471 49755 38477
rect 46400 38440 49648 38468
rect 38565 38403 38623 38409
rect 38565 38369 38577 38403
rect 38611 38400 38623 38403
rect 38654 38400 38660 38412
rect 38611 38372 38660 38400
rect 38611 38369 38623 38372
rect 38565 38363 38623 38369
rect 38654 38360 38660 38372
rect 38712 38360 38718 38412
rect 40126 38400 40132 38412
rect 39132 38372 40132 38400
rect 37918 38332 37924 38344
rect 37879 38304 37924 38332
rect 37918 38292 37924 38304
rect 37976 38292 37982 38344
rect 38102 38292 38108 38344
rect 38160 38332 38166 38344
rect 39132 38341 39160 38372
rect 40126 38360 40132 38372
rect 40184 38400 40190 38412
rect 41874 38400 41880 38412
rect 40184 38372 41880 38400
rect 40184 38360 40190 38372
rect 39117 38335 39175 38341
rect 39117 38332 39129 38335
rect 38160 38304 39129 38332
rect 38160 38292 38166 38304
rect 39117 38301 39129 38304
rect 39163 38301 39175 38335
rect 39117 38295 39175 38301
rect 39301 38335 39359 38341
rect 39301 38301 39313 38335
rect 39347 38332 39359 38335
rect 39482 38332 39488 38344
rect 39347 38304 39488 38332
rect 39347 38301 39359 38304
rect 39301 38295 39359 38301
rect 39482 38292 39488 38304
rect 39540 38292 39546 38344
rect 39758 38292 39764 38344
rect 39816 38332 39822 38344
rect 40512 38341 40540 38372
rect 41874 38360 41880 38372
rect 41932 38360 41938 38412
rect 42518 38360 42524 38412
rect 42576 38400 42582 38412
rect 43441 38403 43499 38409
rect 43441 38400 43453 38403
rect 42576 38372 43453 38400
rect 42576 38360 42582 38372
rect 43441 38369 43453 38372
rect 43487 38369 43499 38403
rect 45738 38400 45744 38412
rect 45699 38372 45744 38400
rect 43441 38363 43499 38369
rect 45738 38360 45744 38372
rect 45796 38360 45802 38412
rect 46400 38409 46428 38440
rect 46385 38403 46443 38409
rect 46385 38369 46397 38403
rect 46431 38369 46443 38403
rect 46385 38363 46443 38369
rect 47210 38360 47216 38412
rect 47268 38400 47274 38412
rect 49050 38400 49056 38412
rect 47268 38372 49056 38400
rect 47268 38360 47274 38372
rect 49050 38360 49056 38372
rect 49108 38360 49114 38412
rect 49234 38400 49240 38412
rect 49195 38372 49240 38400
rect 49234 38360 49240 38372
rect 49292 38360 49298 38412
rect 49620 38400 49648 38440
rect 49697 38437 49709 38471
rect 49743 38468 49755 38471
rect 51166 38468 51172 38480
rect 49743 38440 51172 38468
rect 49743 38437 49755 38440
rect 49697 38431 49755 38437
rect 51166 38428 51172 38440
rect 51224 38428 51230 38480
rect 53834 38428 53840 38480
rect 53892 38468 53898 38480
rect 54573 38471 54631 38477
rect 54573 38468 54585 38471
rect 53892 38440 54585 38468
rect 53892 38428 53898 38440
rect 54220 38412 54248 38440
rect 54573 38437 54585 38440
rect 54619 38468 54631 38471
rect 54846 38468 54852 38480
rect 54619 38440 54852 38468
rect 54619 38437 54631 38440
rect 54573 38431 54631 38437
rect 54846 38428 54852 38440
rect 54904 38428 54910 38480
rect 52825 38403 52883 38409
rect 49620 38372 51074 38400
rect 40405 38335 40463 38341
rect 40405 38332 40417 38335
rect 39816 38304 40417 38332
rect 39816 38292 39822 38304
rect 40405 38301 40417 38304
rect 40451 38301 40463 38335
rect 40405 38295 40463 38301
rect 40498 38335 40556 38341
rect 40498 38301 40510 38335
rect 40544 38301 40556 38335
rect 40678 38332 40684 38344
rect 40639 38304 40684 38332
rect 40498 38295 40556 38301
rect 40678 38292 40684 38304
rect 40736 38292 40742 38344
rect 40954 38341 40960 38344
rect 40911 38335 40960 38341
rect 40911 38301 40923 38335
rect 40957 38301 40960 38335
rect 40911 38295 40960 38301
rect 40954 38292 40960 38295
rect 41012 38292 41018 38344
rect 43530 38332 43536 38344
rect 43491 38304 43536 38332
rect 43530 38292 43536 38304
rect 43588 38292 43594 38344
rect 45554 38332 45560 38344
rect 45515 38304 45560 38332
rect 45554 38292 45560 38304
rect 45612 38292 45618 38344
rect 46934 38292 46940 38344
rect 46992 38332 46998 38344
rect 47397 38335 47455 38341
rect 47397 38332 47409 38335
rect 46992 38304 47409 38332
rect 46992 38292 46998 38304
rect 47397 38301 47409 38304
rect 47443 38332 47455 38335
rect 47857 38335 47915 38341
rect 47857 38332 47869 38335
rect 47443 38304 47869 38332
rect 47443 38301 47455 38304
rect 47397 38295 47455 38301
rect 47857 38301 47869 38304
rect 47903 38301 47915 38335
rect 47857 38295 47915 38301
rect 49329 38335 49387 38341
rect 49329 38301 49341 38335
rect 49375 38332 49387 38335
rect 49418 38332 49424 38344
rect 49375 38304 49424 38332
rect 49375 38301 49387 38304
rect 49329 38295 49387 38301
rect 49418 38292 49424 38304
rect 49476 38292 49482 38344
rect 50338 38332 50344 38344
rect 50299 38304 50344 38332
rect 50338 38292 50344 38304
rect 50396 38292 50402 38344
rect 50430 38292 50436 38344
rect 50488 38332 50494 38344
rect 50488 38304 50533 38332
rect 50488 38292 50494 38304
rect 50798 38292 50804 38344
rect 50856 38341 50862 38344
rect 50856 38332 50864 38341
rect 51046 38332 51074 38372
rect 52825 38369 52837 38403
rect 52871 38400 52883 38403
rect 53006 38400 53012 38412
rect 52871 38372 53012 38400
rect 52871 38369 52883 38372
rect 52825 38363 52883 38369
rect 53006 38360 53012 38372
rect 53064 38360 53070 38412
rect 53558 38360 53564 38412
rect 53616 38400 53622 38412
rect 54113 38403 54171 38409
rect 54113 38400 54125 38403
rect 53616 38372 54125 38400
rect 53616 38360 53622 38372
rect 54113 38369 54125 38372
rect 54159 38369 54171 38403
rect 54113 38363 54171 38369
rect 54202 38360 54208 38412
rect 54260 38360 54266 38412
rect 55214 38360 55220 38412
rect 55272 38400 55278 38412
rect 55585 38403 55643 38409
rect 55585 38400 55597 38403
rect 55272 38372 55597 38400
rect 55272 38360 55278 38372
rect 55585 38369 55597 38372
rect 55631 38369 55643 38403
rect 55585 38363 55643 38369
rect 52733 38335 52791 38341
rect 52733 38332 52745 38335
rect 50856 38304 50901 38332
rect 51046 38304 52745 38332
rect 50856 38295 50864 38304
rect 52733 38301 52745 38304
rect 52779 38332 52791 38335
rect 53190 38332 53196 38344
rect 52779 38304 53196 38332
rect 52779 38301 52791 38304
rect 52733 38295 52791 38301
rect 50856 38292 50862 38295
rect 53190 38292 53196 38304
rect 53248 38292 53254 38344
rect 53837 38335 53895 38341
rect 53837 38301 53849 38335
rect 53883 38332 53895 38335
rect 54018 38332 54024 38344
rect 53883 38304 54024 38332
rect 53883 38301 53895 38304
rect 53837 38295 53895 38301
rect 40218 38264 40224 38276
rect 37752 38236 40224 38264
rect 36219 38233 36231 38236
rect 36173 38227 36231 38233
rect 31846 38196 31852 38208
rect 30800 38168 31852 38196
rect 30800 38156 30806 38168
rect 31846 38156 31852 38168
rect 31904 38156 31910 38208
rect 35066 38156 35072 38208
rect 35124 38196 35130 38208
rect 36188 38196 36216 38227
rect 40218 38224 40224 38236
rect 40276 38224 40282 38276
rect 40773 38267 40831 38273
rect 40773 38233 40785 38267
rect 40819 38233 40831 38267
rect 40773 38227 40831 38233
rect 41877 38267 41935 38273
rect 41877 38233 41889 38267
rect 41923 38264 41935 38267
rect 42334 38264 42340 38276
rect 41923 38236 42340 38264
rect 41923 38233 41935 38236
rect 41877 38227 41935 38233
rect 36722 38196 36728 38208
rect 35124 38168 36216 38196
rect 36683 38168 36728 38196
rect 35124 38156 35130 38168
rect 36722 38156 36728 38168
rect 36780 38196 36786 38208
rect 37826 38196 37832 38208
rect 36780 38168 37832 38196
rect 36780 38156 36786 38168
rect 37826 38156 37832 38168
rect 37884 38156 37890 38208
rect 39485 38199 39543 38205
rect 39485 38165 39497 38199
rect 39531 38196 39543 38199
rect 39574 38196 39580 38208
rect 39531 38168 39580 38196
rect 39531 38165 39543 38168
rect 39485 38159 39543 38165
rect 39574 38156 39580 38168
rect 39632 38156 39638 38208
rect 40402 38156 40408 38208
rect 40460 38196 40466 38208
rect 40788 38196 40816 38227
rect 42334 38224 42340 38236
rect 42392 38224 42398 38276
rect 42426 38224 42432 38276
rect 42484 38264 42490 38276
rect 42521 38267 42579 38273
rect 42521 38264 42533 38267
rect 42484 38236 42533 38264
rect 42484 38224 42490 38236
rect 42521 38233 42533 38236
rect 42567 38233 42579 38267
rect 42521 38227 42579 38233
rect 42794 38224 42800 38276
rect 42852 38264 42858 38276
rect 42889 38267 42947 38273
rect 42889 38264 42901 38267
rect 42852 38236 42901 38264
rect 42852 38224 42858 38236
rect 42889 38233 42901 38236
rect 42935 38233 42947 38267
rect 42889 38227 42947 38233
rect 47762 38224 47768 38276
rect 47820 38264 47826 38276
rect 48133 38267 48191 38273
rect 48133 38264 48145 38267
rect 47820 38236 48145 38264
rect 47820 38224 47826 38236
rect 48133 38233 48145 38236
rect 48179 38233 48191 38267
rect 48133 38227 48191 38233
rect 50617 38267 50675 38273
rect 50617 38233 50629 38267
rect 50663 38233 50675 38267
rect 50617 38227 50675 38233
rect 40460 38168 40816 38196
rect 41785 38199 41843 38205
rect 40460 38156 40466 38168
rect 41785 38165 41797 38199
rect 41831 38196 41843 38199
rect 42150 38196 42156 38208
rect 41831 38168 42156 38196
rect 41831 38165 41843 38168
rect 41785 38159 41843 38165
rect 42150 38156 42156 38168
rect 42208 38196 42214 38208
rect 45646 38196 45652 38208
rect 42208 38168 45652 38196
rect 42208 38156 42214 38168
rect 45646 38156 45652 38168
rect 45704 38196 45710 38208
rect 47670 38196 47676 38208
rect 45704 38168 47676 38196
rect 45704 38156 45710 38168
rect 47670 38156 47676 38168
rect 47728 38196 47734 38208
rect 47949 38199 48007 38205
rect 47949 38196 47961 38199
rect 47728 38168 47961 38196
rect 47728 38156 47734 38168
rect 47949 38165 47961 38168
rect 47995 38165 48007 38199
rect 48682 38196 48688 38208
rect 48643 38168 48688 38196
rect 47949 38159 48007 38165
rect 48682 38156 48688 38168
rect 48740 38156 48746 38208
rect 50632 38196 50660 38227
rect 50706 38224 50712 38276
rect 50764 38264 50770 38276
rect 50764 38236 50809 38264
rect 50764 38224 50770 38236
rect 50890 38224 50896 38276
rect 50948 38264 50954 38276
rect 51445 38267 51503 38273
rect 51445 38264 51457 38267
rect 50948 38236 51457 38264
rect 50948 38224 50954 38236
rect 51445 38233 51457 38236
rect 51491 38233 51503 38267
rect 51445 38227 51503 38233
rect 52362 38224 52368 38276
rect 52420 38264 52426 38276
rect 53852 38264 53880 38295
rect 54018 38292 54024 38304
rect 54076 38292 54082 38344
rect 55674 38332 55680 38344
rect 55635 38304 55680 38332
rect 55674 38292 55680 38304
rect 55732 38292 55738 38344
rect 52420 38236 53880 38264
rect 52420 38224 52426 38236
rect 51994 38196 52000 38208
rect 50632 38168 52000 38196
rect 51994 38156 52000 38168
rect 52052 38156 52058 38208
rect 53101 38199 53159 38205
rect 53101 38165 53113 38199
rect 53147 38196 53159 38199
rect 54478 38196 54484 38208
rect 53147 38168 54484 38196
rect 53147 38165 53159 38168
rect 53101 38159 53159 38165
rect 54478 38156 54484 38168
rect 54536 38156 54542 38208
rect 56042 38196 56048 38208
rect 56003 38168 56048 38196
rect 56042 38156 56048 38168
rect 56100 38156 56106 38208
rect 1104 38106 58880 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 35594 38106
rect 35646 38054 35658 38106
rect 35710 38054 35722 38106
rect 35774 38054 35786 38106
rect 35838 38054 35850 38106
rect 35902 38054 58880 38106
rect 1104 38032 58880 38054
rect 29270 37992 29276 38004
rect 29231 37964 29276 37992
rect 29270 37952 29276 37964
rect 29328 37952 29334 38004
rect 31478 37952 31484 38004
rect 31536 37992 31542 38004
rect 31665 37995 31723 38001
rect 31665 37992 31677 37995
rect 31536 37964 31677 37992
rect 31536 37952 31542 37964
rect 31665 37961 31677 37964
rect 31711 37961 31723 37995
rect 31665 37955 31723 37961
rect 32769 37995 32827 38001
rect 32769 37961 32781 37995
rect 32815 37992 32827 37995
rect 33042 37992 33048 38004
rect 32815 37964 33048 37992
rect 32815 37961 32827 37964
rect 32769 37955 32827 37961
rect 33042 37952 33048 37964
rect 33100 37952 33106 38004
rect 33413 37995 33471 38001
rect 33413 37961 33425 37995
rect 33459 37961 33471 37995
rect 33413 37955 33471 37961
rect 34425 37995 34483 38001
rect 34425 37961 34437 37995
rect 34471 37992 34483 37995
rect 34790 37992 34796 38004
rect 34471 37964 34796 37992
rect 34471 37961 34483 37964
rect 34425 37955 34483 37961
rect 30558 37924 30564 37936
rect 30116 37896 30564 37924
rect 29178 37856 29184 37868
rect 29139 37828 29184 37856
rect 29178 37816 29184 37828
rect 29236 37816 29242 37868
rect 30116 37865 30144 37896
rect 30558 37884 30564 37896
rect 30616 37924 30622 37936
rect 31938 37924 31944 37936
rect 30616 37896 31944 37924
rect 30616 37884 30622 37896
rect 31938 37884 31944 37896
rect 31996 37884 32002 37936
rect 32490 37924 32496 37936
rect 32403 37896 32496 37924
rect 32490 37884 32496 37896
rect 32548 37924 32554 37936
rect 33428 37924 33456 37955
rect 34790 37952 34796 37964
rect 34848 37952 34854 38004
rect 38930 37992 38936 38004
rect 38626 37964 38936 37992
rect 32548 37896 33456 37924
rect 32548 37884 32554 37896
rect 33502 37884 33508 37936
rect 33560 37933 33566 37936
rect 33560 37927 33623 37933
rect 33560 37893 33577 37927
rect 33611 37893 33623 37927
rect 33560 37887 33623 37893
rect 33560 37884 33566 37887
rect 33686 37884 33692 37936
rect 33744 37924 33750 37936
rect 33781 37927 33839 37933
rect 33781 37924 33793 37927
rect 33744 37896 33793 37924
rect 33744 37884 33750 37896
rect 33781 37893 33793 37896
rect 33827 37893 33839 37927
rect 35526 37924 35532 37936
rect 33781 37887 33839 37893
rect 34808 37896 35532 37924
rect 30101 37859 30159 37865
rect 30101 37825 30113 37859
rect 30147 37825 30159 37859
rect 30101 37819 30159 37825
rect 30374 37816 30380 37868
rect 30432 37856 30438 37868
rect 30469 37859 30527 37865
rect 30469 37856 30481 37859
rect 30432 37828 30481 37856
rect 30432 37816 30438 37828
rect 30469 37825 30481 37828
rect 30515 37825 30527 37859
rect 30926 37856 30932 37868
rect 30887 37828 30932 37856
rect 30469 37819 30527 37825
rect 30190 37788 30196 37800
rect 30151 37760 30196 37788
rect 30190 37748 30196 37760
rect 30248 37748 30254 37800
rect 30484 37788 30512 37819
rect 30926 37816 30932 37828
rect 30984 37816 30990 37868
rect 31202 37816 31208 37868
rect 31260 37856 31266 37868
rect 31481 37859 31539 37865
rect 31481 37856 31493 37859
rect 31260 37828 31493 37856
rect 31260 37816 31266 37828
rect 31481 37825 31493 37828
rect 31527 37825 31539 37859
rect 31481 37819 31539 37825
rect 31570 37816 31576 37868
rect 31628 37856 31634 37868
rect 32508 37856 32536 37884
rect 34808 37865 34836 37896
rect 35526 37884 35532 37896
rect 35584 37924 35590 37936
rect 35986 37924 35992 37936
rect 35584 37896 35894 37924
rect 35947 37896 35992 37924
rect 35584 37884 35590 37896
rect 31628 37828 32536 37856
rect 34609 37859 34667 37865
rect 31628 37816 31634 37828
rect 34609 37825 34621 37859
rect 34655 37825 34667 37859
rect 34609 37819 34667 37825
rect 34793 37859 34851 37865
rect 34793 37825 34805 37859
rect 34839 37825 34851 37859
rect 34793 37819 34851 37825
rect 34885 37859 34943 37865
rect 34885 37825 34897 37859
rect 34931 37825 34943 37859
rect 34885 37819 34943 37825
rect 30834 37788 30840 37800
rect 30484 37760 30840 37788
rect 30834 37748 30840 37760
rect 30892 37748 30898 37800
rect 28721 37655 28779 37661
rect 28721 37621 28733 37655
rect 28767 37652 28779 37655
rect 29270 37652 29276 37664
rect 28767 37624 29276 37652
rect 28767 37621 28779 37624
rect 28721 37615 28779 37621
rect 29270 37612 29276 37624
rect 29328 37612 29334 37664
rect 33597 37655 33655 37661
rect 33597 37621 33609 37655
rect 33643 37652 33655 37655
rect 33778 37652 33784 37664
rect 33643 37624 33784 37652
rect 33643 37621 33655 37624
rect 33597 37615 33655 37621
rect 33778 37612 33784 37624
rect 33836 37612 33842 37664
rect 34624 37652 34652 37819
rect 34900 37788 34928 37819
rect 34974 37816 34980 37868
rect 35032 37856 35038 37868
rect 35345 37859 35403 37865
rect 35345 37856 35357 37859
rect 35032 37828 35357 37856
rect 35032 37816 35038 37828
rect 35345 37825 35357 37828
rect 35391 37825 35403 37859
rect 35345 37819 35403 37825
rect 35434 37816 35440 37868
rect 35492 37856 35498 37868
rect 35621 37859 35679 37865
rect 35621 37856 35633 37859
rect 35492 37828 35633 37856
rect 35492 37816 35498 37828
rect 35621 37825 35633 37828
rect 35667 37825 35679 37859
rect 35866 37856 35894 37896
rect 35986 37884 35992 37896
rect 36044 37884 36050 37936
rect 38626 37924 38654 37964
rect 38930 37952 38936 37964
rect 38988 37952 38994 38004
rect 39482 37952 39488 38004
rect 39540 37952 39546 38004
rect 39758 37992 39764 38004
rect 39719 37964 39764 37992
rect 39758 37952 39764 37964
rect 39816 37952 39822 38004
rect 40770 37952 40776 38004
rect 40828 37992 40834 38004
rect 41690 37992 41696 38004
rect 40828 37964 41696 37992
rect 40828 37952 40834 37964
rect 41690 37952 41696 37964
rect 41748 37952 41754 38004
rect 41874 37952 41880 38004
rect 41932 37992 41938 38004
rect 42242 37992 42248 38004
rect 41932 37964 42248 37992
rect 41932 37952 41938 37964
rect 42242 37952 42248 37964
rect 42300 37992 42306 38004
rect 42300 37964 43024 37992
rect 42300 37952 42306 37964
rect 36280 37896 38654 37924
rect 39500 37924 39528 37952
rect 39500 37896 39804 37924
rect 36280 37856 36308 37896
rect 35866 37828 36308 37856
rect 35621 37819 35679 37825
rect 36354 37816 36360 37868
rect 36412 37856 36418 37868
rect 36449 37859 36507 37865
rect 36449 37856 36461 37859
rect 36412 37828 36461 37856
rect 36412 37816 36418 37828
rect 36449 37825 36461 37828
rect 36495 37825 36507 37859
rect 36630 37856 36636 37868
rect 36591 37828 36636 37856
rect 36449 37819 36507 37825
rect 36630 37816 36636 37828
rect 36688 37816 36694 37868
rect 37476 37865 37504 37896
rect 37461 37859 37519 37865
rect 37461 37825 37473 37859
rect 37507 37825 37519 37859
rect 37461 37819 37519 37825
rect 37645 37859 37703 37865
rect 37645 37825 37657 37859
rect 37691 37825 37703 37859
rect 37645 37819 37703 37825
rect 35805 37791 35863 37797
rect 35805 37788 35817 37791
rect 34900 37760 35817 37788
rect 35805 37757 35817 37760
rect 35851 37788 35863 37791
rect 36541 37791 36599 37797
rect 36541 37788 36553 37791
rect 35851 37760 36553 37788
rect 35851 37757 35863 37760
rect 35805 37751 35863 37757
rect 36541 37757 36553 37760
rect 36587 37788 36599 37791
rect 37660 37788 37688 37819
rect 37826 37816 37832 37868
rect 37884 37856 37890 37868
rect 37921 37859 37979 37865
rect 37921 37856 37933 37859
rect 37884 37828 37933 37856
rect 37884 37816 37890 37828
rect 37921 37825 37933 37828
rect 37967 37825 37979 37859
rect 39482 37856 39488 37868
rect 39443 37828 39488 37856
rect 37921 37819 37979 37825
rect 39482 37816 39488 37828
rect 39540 37816 39546 37868
rect 39577 37859 39635 37865
rect 39577 37825 39589 37859
rect 39623 37856 39635 37859
rect 39666 37856 39672 37868
rect 39623 37828 39672 37856
rect 39623 37825 39635 37828
rect 39577 37819 39635 37825
rect 39666 37816 39672 37828
rect 39724 37816 39730 37868
rect 39776 37797 39804 37896
rect 40218 37884 40224 37936
rect 40276 37924 40282 37936
rect 40313 37927 40371 37933
rect 40313 37924 40325 37927
rect 40276 37896 40325 37924
rect 40276 37884 40282 37896
rect 40313 37893 40325 37896
rect 40359 37893 40371 37927
rect 42886 37924 42892 37936
rect 40313 37887 40371 37893
rect 41248 37896 42748 37924
rect 42847 37896 42892 37924
rect 36587 37760 37688 37788
rect 39761 37791 39819 37797
rect 36587 37757 36599 37760
rect 36541 37751 36599 37757
rect 39761 37757 39773 37791
rect 39807 37757 39819 37791
rect 40328 37788 40356 37887
rect 40402 37816 40408 37868
rect 40460 37856 40466 37868
rect 41248 37865 41276 37896
rect 42720 37868 42748 37896
rect 42886 37884 42892 37896
rect 42944 37884 42950 37936
rect 42996 37933 43024 37964
rect 51902 37952 51908 38004
rect 51960 37992 51966 38004
rect 52273 37995 52331 38001
rect 52273 37992 52285 37995
rect 51960 37964 52285 37992
rect 51960 37952 51966 37964
rect 52273 37961 52285 37964
rect 52319 37992 52331 37995
rect 52362 37992 52368 38004
rect 52319 37964 52368 37992
rect 52319 37961 52331 37964
rect 52273 37955 52331 37961
rect 52362 37952 52368 37964
rect 52420 37952 52426 38004
rect 54110 37952 54116 38004
rect 54168 37992 54174 38004
rect 54481 37995 54539 38001
rect 54481 37992 54493 37995
rect 54168 37964 54493 37992
rect 54168 37952 54174 37964
rect 54481 37961 54493 37964
rect 54527 37961 54539 37995
rect 54481 37955 54539 37961
rect 54846 37952 54852 38004
rect 54904 37992 54910 38004
rect 55033 37995 55091 38001
rect 55033 37992 55045 37995
rect 54904 37964 55045 37992
rect 54904 37952 54910 37964
rect 55033 37961 55045 37964
rect 55079 37961 55091 37995
rect 55033 37955 55091 37961
rect 42981 37927 43039 37933
rect 42981 37893 42993 37927
rect 43027 37893 43039 37927
rect 43806 37924 43812 37936
rect 43719 37896 43812 37924
rect 42981 37887 43039 37893
rect 43806 37884 43812 37896
rect 43864 37924 43870 37936
rect 45278 37924 45284 37936
rect 43864 37896 45284 37924
rect 43864 37884 43870 37896
rect 45278 37884 45284 37896
rect 45336 37884 45342 37936
rect 47029 37927 47087 37933
rect 47029 37924 47041 37927
rect 45572 37896 47041 37924
rect 41233 37859 41291 37865
rect 41233 37856 41245 37859
rect 40460 37828 41245 37856
rect 40460 37816 40466 37828
rect 41233 37825 41245 37828
rect 41279 37825 41291 37859
rect 42610 37856 42616 37868
rect 42571 37828 42616 37856
rect 41233 37819 41291 37825
rect 42610 37816 42616 37828
rect 42668 37816 42674 37868
rect 42702 37816 42708 37868
rect 42760 37856 42766 37868
rect 42760 37828 42805 37856
rect 42760 37816 42766 37828
rect 43070 37816 43076 37868
rect 43128 37865 43134 37868
rect 43128 37856 43136 37865
rect 44821 37859 44879 37865
rect 44821 37856 44833 37859
rect 43128 37828 43173 37856
rect 43272 37828 44833 37856
rect 43128 37819 43136 37828
rect 43128 37816 43134 37819
rect 42058 37788 42064 37800
rect 40328 37760 42064 37788
rect 39761 37751 39819 37757
rect 42058 37748 42064 37760
rect 42116 37748 42122 37800
rect 42518 37748 42524 37800
rect 42576 37788 42582 37800
rect 43272 37788 43300 37828
rect 44821 37825 44833 37828
rect 44867 37825 44879 37859
rect 44821 37819 44879 37825
rect 42576 37760 43300 37788
rect 42576 37748 42582 37760
rect 43714 37748 43720 37800
rect 43772 37788 43778 37800
rect 44729 37791 44787 37797
rect 44729 37788 44741 37791
rect 43772 37760 44741 37788
rect 43772 37748 43778 37760
rect 44729 37757 44741 37760
rect 44775 37757 44787 37791
rect 44729 37751 44787 37757
rect 38105 37723 38163 37729
rect 38105 37689 38117 37723
rect 38151 37720 38163 37723
rect 39942 37720 39948 37732
rect 38151 37692 39948 37720
rect 38151 37689 38163 37692
rect 38105 37683 38163 37689
rect 39942 37680 39948 37692
rect 40000 37680 40006 37732
rect 41690 37680 41696 37732
rect 41748 37720 41754 37732
rect 45572 37720 45600 37896
rect 47029 37893 47041 37896
rect 47075 37924 47087 37927
rect 48314 37924 48320 37936
rect 47075 37896 48320 37924
rect 47075 37893 47087 37896
rect 47029 37887 47087 37893
rect 48314 37884 48320 37896
rect 48372 37924 48378 37936
rect 48501 37927 48559 37933
rect 48501 37924 48513 37927
rect 48372 37896 48513 37924
rect 48372 37884 48378 37896
rect 48501 37893 48513 37896
rect 48547 37924 48559 37927
rect 48682 37924 48688 37936
rect 48547 37896 48688 37924
rect 48547 37893 48559 37896
rect 48501 37887 48559 37893
rect 48682 37884 48688 37896
rect 48740 37924 48746 37936
rect 49237 37927 49295 37933
rect 49237 37924 49249 37927
rect 48740 37896 49249 37924
rect 48740 37884 48746 37896
rect 49237 37893 49249 37896
rect 49283 37924 49295 37927
rect 49326 37924 49332 37936
rect 49283 37896 49332 37924
rect 49283 37893 49295 37896
rect 49237 37887 49295 37893
rect 49326 37884 49332 37896
rect 49384 37884 49390 37936
rect 54021 37927 54079 37933
rect 54021 37893 54033 37927
rect 54067 37924 54079 37927
rect 56134 37924 56140 37936
rect 54067 37896 56140 37924
rect 54067 37893 54079 37896
rect 54021 37887 54079 37893
rect 56134 37884 56140 37896
rect 56192 37884 56198 37936
rect 46106 37816 46112 37868
rect 46164 37856 46170 37868
rect 46293 37859 46351 37865
rect 46293 37856 46305 37859
rect 46164 37828 46305 37856
rect 46164 37816 46170 37828
rect 46293 37825 46305 37828
rect 46339 37825 46351 37859
rect 46293 37819 46351 37825
rect 46477 37859 46535 37865
rect 46477 37825 46489 37859
rect 46523 37825 46535 37859
rect 46934 37856 46940 37868
rect 46895 37828 46940 37856
rect 46477 37819 46535 37825
rect 45649 37791 45707 37797
rect 45649 37757 45661 37791
rect 45695 37757 45707 37791
rect 45649 37751 45707 37757
rect 41748 37692 45600 37720
rect 45664 37720 45692 37751
rect 46014 37748 46020 37800
rect 46072 37788 46078 37800
rect 46492 37788 46520 37819
rect 46934 37816 46940 37828
rect 46992 37816 46998 37868
rect 47213 37859 47271 37865
rect 47213 37825 47225 37859
rect 47259 37856 47271 37859
rect 47762 37856 47768 37868
rect 47259 37828 47768 37856
rect 47259 37825 47271 37828
rect 47213 37819 47271 37825
rect 47762 37816 47768 37828
rect 47820 37816 47826 37868
rect 48133 37859 48191 37865
rect 48133 37825 48145 37859
rect 48179 37825 48191 37859
rect 48133 37819 48191 37825
rect 48148 37788 48176 37819
rect 48222 37816 48228 37868
rect 48280 37856 48286 37868
rect 48280 37828 48325 37856
rect 48280 37816 48286 37828
rect 48406 37816 48412 37868
rect 48464 37856 48470 37868
rect 48464 37828 48509 37856
rect 48464 37816 48470 37828
rect 48590 37816 48596 37868
rect 48648 37865 48654 37868
rect 48648 37856 48656 37865
rect 50893 37859 50951 37865
rect 50893 37856 50905 37859
rect 48648 37828 48693 37856
rect 48792 37828 50905 37856
rect 48648 37819 48656 37828
rect 48648 37816 48654 37819
rect 46072 37760 46520 37788
rect 47228 37760 48176 37788
rect 46072 37748 46078 37760
rect 47228 37729 47256 37760
rect 48792 37729 48820 37828
rect 50893 37825 50905 37828
rect 50939 37825 50951 37859
rect 53190 37856 53196 37868
rect 53151 37828 53196 37856
rect 50893 37819 50951 37825
rect 53190 37816 53196 37828
rect 53248 37816 53254 37868
rect 55950 37856 55956 37868
rect 55911 37828 55956 37856
rect 55950 37816 55956 37828
rect 56008 37816 56014 37868
rect 56318 37816 56324 37868
rect 56376 37856 56382 37868
rect 56965 37859 57023 37865
rect 56965 37856 56977 37859
rect 56376 37828 56977 37856
rect 56376 37816 56382 37828
rect 56965 37825 56977 37828
rect 57011 37825 57023 37859
rect 56965 37819 57023 37825
rect 50798 37788 50804 37800
rect 49160 37760 50804 37788
rect 47213 37723 47271 37729
rect 45664 37692 47164 37720
rect 41748 37680 41754 37692
rect 35342 37652 35348 37664
rect 34624 37624 35348 37652
rect 35342 37612 35348 37624
rect 35400 37612 35406 37664
rect 37550 37612 37556 37664
rect 37608 37652 37614 37664
rect 38657 37655 38715 37661
rect 38657 37652 38669 37655
rect 37608 37624 38669 37652
rect 37608 37612 37614 37624
rect 38657 37621 38669 37624
rect 38703 37621 38715 37655
rect 38657 37615 38715 37621
rect 39482 37612 39488 37664
rect 39540 37652 39546 37664
rect 40402 37652 40408 37664
rect 39540 37624 40408 37652
rect 39540 37612 39546 37624
rect 40402 37612 40408 37624
rect 40460 37612 40466 37664
rect 40589 37655 40647 37661
rect 40589 37621 40601 37655
rect 40635 37652 40647 37655
rect 40770 37652 40776 37664
rect 40635 37624 40776 37652
rect 40635 37621 40647 37624
rect 40589 37615 40647 37621
rect 40770 37612 40776 37624
rect 40828 37612 40834 37664
rect 41509 37655 41567 37661
rect 41509 37621 41521 37655
rect 41555 37652 41567 37655
rect 41966 37652 41972 37664
rect 41555 37624 41972 37652
rect 41555 37621 41567 37624
rect 41509 37615 41567 37621
rect 41966 37612 41972 37624
rect 42024 37612 42030 37664
rect 43257 37655 43315 37661
rect 43257 37621 43269 37655
rect 43303 37652 43315 37655
rect 43346 37652 43352 37664
rect 43303 37624 43352 37652
rect 43303 37621 43315 37624
rect 43257 37615 43315 37621
rect 43346 37612 43352 37624
rect 43404 37612 43410 37664
rect 46474 37652 46480 37664
rect 46435 37624 46480 37652
rect 46474 37612 46480 37624
rect 46532 37612 46538 37664
rect 47136 37652 47164 37692
rect 47213 37689 47225 37723
rect 47259 37689 47271 37723
rect 47213 37683 47271 37689
rect 48777 37723 48835 37729
rect 48777 37689 48789 37723
rect 48823 37689 48835 37723
rect 48777 37683 48835 37689
rect 49160 37652 49188 37760
rect 50798 37748 50804 37760
rect 50856 37748 50862 37800
rect 51261 37791 51319 37797
rect 51261 37757 51273 37791
rect 51307 37788 51319 37791
rect 53101 37791 53159 37797
rect 53101 37788 53113 37791
rect 51307 37760 53113 37788
rect 51307 37757 51319 37760
rect 51261 37751 51319 37757
rect 53101 37757 53113 37760
rect 53147 37757 53159 37791
rect 53101 37751 53159 37757
rect 54478 37748 54484 37800
rect 54536 37788 54542 37800
rect 55858 37788 55864 37800
rect 54536 37760 55864 37788
rect 54536 37748 54542 37760
rect 55858 37748 55864 37760
rect 55916 37748 55922 37800
rect 56042 37748 56048 37800
rect 56100 37788 56106 37800
rect 56873 37791 56931 37797
rect 56873 37788 56885 37791
rect 56100 37760 56885 37788
rect 56100 37748 56106 37760
rect 56873 37757 56885 37760
rect 56919 37757 56931 37791
rect 56873 37751 56931 37757
rect 56321 37723 56379 37729
rect 56321 37689 56333 37723
rect 56367 37720 56379 37723
rect 57698 37720 57704 37732
rect 56367 37692 57704 37720
rect 56367 37689 56379 37692
rect 56321 37683 56379 37689
rect 57698 37680 57704 37692
rect 57756 37680 57762 37732
rect 49786 37652 49792 37664
rect 47136 37624 49188 37652
rect 49747 37624 49792 37652
rect 49786 37612 49792 37624
rect 49844 37652 49850 37664
rect 50430 37652 50436 37664
rect 49844 37624 50436 37652
rect 49844 37612 49850 37624
rect 50430 37612 50436 37624
rect 50488 37652 50494 37664
rect 50890 37652 50896 37664
rect 50488 37624 50896 37652
rect 50488 37612 50494 37624
rect 50890 37612 50896 37624
rect 50948 37612 50954 37664
rect 57238 37652 57244 37664
rect 57199 37624 57244 37652
rect 57238 37612 57244 37624
rect 57296 37612 57302 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 29181 37451 29239 37457
rect 29181 37417 29193 37451
rect 29227 37448 29239 37451
rect 30650 37448 30656 37460
rect 29227 37420 30656 37448
rect 29227 37417 29239 37420
rect 29181 37411 29239 37417
rect 30650 37408 30656 37420
rect 30708 37408 30714 37460
rect 32306 37448 32312 37460
rect 32267 37420 32312 37448
rect 32306 37408 32312 37420
rect 32364 37408 32370 37460
rect 32674 37408 32680 37460
rect 32732 37408 32738 37460
rect 32766 37408 32772 37460
rect 32824 37448 32830 37460
rect 34885 37451 34943 37457
rect 34885 37448 34897 37451
rect 32824 37420 34897 37448
rect 32824 37408 32830 37420
rect 34885 37417 34897 37420
rect 34931 37417 34943 37451
rect 34885 37411 34943 37417
rect 37369 37451 37427 37457
rect 37369 37417 37381 37451
rect 37415 37448 37427 37451
rect 37458 37448 37464 37460
rect 37415 37420 37464 37448
rect 37415 37417 37427 37420
rect 37369 37411 37427 37417
rect 37458 37408 37464 37420
rect 37516 37448 37522 37460
rect 37642 37448 37648 37460
rect 37516 37420 37648 37448
rect 37516 37408 37522 37420
rect 37642 37408 37648 37420
rect 37700 37408 37706 37460
rect 38102 37408 38108 37460
rect 38160 37448 38166 37460
rect 41509 37451 41567 37457
rect 38160 37420 40448 37448
rect 38160 37408 38166 37420
rect 28445 37383 28503 37389
rect 28445 37349 28457 37383
rect 28491 37349 28503 37383
rect 32692 37380 32720 37408
rect 33413 37383 33471 37389
rect 33413 37380 33425 37383
rect 32692 37352 33425 37380
rect 28445 37343 28503 37349
rect 33413 37349 33425 37352
rect 33459 37349 33471 37383
rect 33413 37343 33471 37349
rect 28166 37244 28172 37256
rect 28127 37216 28172 37244
rect 28166 37204 28172 37216
rect 28224 37204 28230 37256
rect 28460 37244 28488 37343
rect 34054 37340 34060 37392
rect 34112 37380 34118 37392
rect 34241 37383 34299 37389
rect 34241 37380 34253 37383
rect 34112 37352 34253 37380
rect 34112 37340 34118 37352
rect 34241 37349 34253 37352
rect 34287 37380 34299 37383
rect 35618 37380 35624 37392
rect 34287 37352 35624 37380
rect 34287 37349 34299 37352
rect 34241 37343 34299 37349
rect 35618 37340 35624 37352
rect 35676 37340 35682 37392
rect 36630 37380 36636 37392
rect 36096 37352 36636 37380
rect 28810 37272 28816 37324
rect 28868 37312 28874 37324
rect 29362 37312 29368 37324
rect 28868 37284 28948 37312
rect 28868 37272 28874 37284
rect 28920 37253 28948 37284
rect 29012 37284 29368 37312
rect 29012 37253 29040 37284
rect 29362 37272 29368 37284
rect 29420 37272 29426 37324
rect 30742 37312 30748 37324
rect 30703 37284 30748 37312
rect 30742 37272 30748 37284
rect 30800 37272 30806 37324
rect 30926 37312 30932 37324
rect 30887 37284 30932 37312
rect 30926 37272 30932 37284
rect 30984 37272 30990 37324
rect 32674 37272 32680 37324
rect 32732 37312 32738 37324
rect 32769 37315 32827 37321
rect 32769 37312 32781 37315
rect 32732 37284 32781 37312
rect 32732 37272 32738 37284
rect 32769 37281 32781 37284
rect 32815 37312 32827 37315
rect 33870 37312 33876 37324
rect 32815 37284 33876 37312
rect 32815 37281 32827 37284
rect 32769 37275 32827 37281
rect 33870 37272 33876 37284
rect 33928 37272 33934 37324
rect 36096 37312 36124 37352
rect 36630 37340 36636 37352
rect 36688 37340 36694 37392
rect 39485 37383 39543 37389
rect 39485 37349 39497 37383
rect 39531 37380 39543 37383
rect 39666 37380 39672 37392
rect 39531 37352 39672 37380
rect 39531 37349 39543 37352
rect 39485 37343 39543 37349
rect 39666 37340 39672 37352
rect 39724 37340 39730 37392
rect 40420 37389 40448 37420
rect 41509 37417 41521 37451
rect 41555 37448 41567 37451
rect 42610 37448 42616 37460
rect 41555 37420 42616 37448
rect 41555 37417 41567 37420
rect 41509 37411 41567 37417
rect 42610 37408 42616 37420
rect 42668 37408 42674 37460
rect 43714 37448 43720 37460
rect 43675 37420 43720 37448
rect 43714 37408 43720 37420
rect 43772 37408 43778 37460
rect 46569 37451 46627 37457
rect 46569 37417 46581 37451
rect 46615 37448 46627 37451
rect 46934 37448 46940 37460
rect 46615 37420 46940 37448
rect 46615 37417 46627 37420
rect 46569 37411 46627 37417
rect 46934 37408 46940 37420
rect 46992 37408 46998 37460
rect 52454 37408 52460 37460
rect 52512 37448 52518 37460
rect 53466 37448 53472 37460
rect 52512 37420 53472 37448
rect 52512 37408 52518 37420
rect 53466 37408 53472 37420
rect 53524 37408 53530 37460
rect 56318 37448 56324 37460
rect 56279 37420 56324 37448
rect 56318 37408 56324 37420
rect 56376 37408 56382 37460
rect 40405 37383 40463 37389
rect 40405 37349 40417 37383
rect 40451 37349 40463 37383
rect 40405 37343 40463 37349
rect 40678 37340 40684 37392
rect 40736 37380 40742 37392
rect 47765 37383 47823 37389
rect 40736 37352 47532 37380
rect 40736 37340 40742 37352
rect 36722 37312 36728 37324
rect 34900 37284 36124 37312
rect 36188 37284 36728 37312
rect 28905 37247 28963 37253
rect 28460 37216 28856 37244
rect 28445 37179 28503 37185
rect 28445 37145 28457 37179
rect 28491 37145 28503 37179
rect 28828 37176 28856 37216
rect 28905 37213 28917 37247
rect 28951 37213 28963 37247
rect 28905 37207 28963 37213
rect 28997 37247 29055 37253
rect 28997 37213 29009 37247
rect 29043 37213 29055 37247
rect 29733 37247 29791 37253
rect 29733 37244 29745 37247
rect 28997 37207 29055 37213
rect 29104 37216 29745 37244
rect 29104 37176 29132 37216
rect 29733 37213 29745 37216
rect 29779 37213 29791 37247
rect 30558 37244 30564 37256
rect 30519 37216 30564 37244
rect 29733 37207 29791 37213
rect 30558 37204 30564 37216
rect 30616 37204 30622 37256
rect 31021 37247 31079 37253
rect 31021 37213 31033 37247
rect 31067 37213 31079 37247
rect 31021 37207 31079 37213
rect 32585 37247 32643 37253
rect 32585 37213 32597 37247
rect 32631 37244 32643 37247
rect 33413 37247 33471 37253
rect 32631 37216 33088 37244
rect 32631 37213 32643 37216
rect 32585 37207 32643 37213
rect 28828 37148 29132 37176
rect 29181 37179 29239 37185
rect 28445 37139 28503 37145
rect 29181 37145 29193 37179
rect 29227 37176 29239 37179
rect 29270 37176 29276 37188
rect 29227 37148 29276 37176
rect 29227 37145 29239 37148
rect 29181 37139 29239 37145
rect 28258 37108 28264 37120
rect 28219 37080 28264 37108
rect 28258 37068 28264 37080
rect 28316 37068 28322 37120
rect 28460 37108 28488 37139
rect 29270 37136 29276 37148
rect 29328 37136 29334 37188
rect 30190 37136 30196 37188
rect 30248 37176 30254 37188
rect 31036 37176 31064 37207
rect 30248 37148 31064 37176
rect 32217 37179 32275 37185
rect 30248 37136 30254 37148
rect 32217 37145 32229 37179
rect 32263 37176 32275 37179
rect 32950 37176 32956 37188
rect 32263 37148 32956 37176
rect 32263 37145 32275 37148
rect 32217 37139 32275 37145
rect 32950 37136 32956 37148
rect 33008 37136 33014 37188
rect 28902 37108 28908 37120
rect 28460 37080 28908 37108
rect 28902 37068 28908 37080
rect 28960 37068 28966 37120
rect 29086 37068 29092 37120
rect 29144 37108 29150 37120
rect 29825 37111 29883 37117
rect 29825 37108 29837 37111
rect 29144 37080 29837 37108
rect 29144 37068 29150 37080
rect 29825 37077 29837 37080
rect 29871 37077 29883 37111
rect 33060 37108 33088 37216
rect 33413 37213 33425 37247
rect 33459 37244 33471 37247
rect 33502 37244 33508 37256
rect 33459 37216 33508 37244
rect 33459 37213 33471 37216
rect 33413 37207 33471 37213
rect 33134 37136 33140 37188
rect 33192 37176 33198 37188
rect 33428 37176 33456 37207
rect 33502 37204 33508 37216
rect 33560 37204 33566 37256
rect 33597 37247 33655 37253
rect 33597 37213 33609 37247
rect 33643 37244 33655 37247
rect 33686 37244 33692 37256
rect 33643 37216 33692 37244
rect 33643 37213 33655 37216
rect 33597 37207 33655 37213
rect 33686 37204 33692 37216
rect 33744 37204 33750 37256
rect 34606 37204 34612 37256
rect 34664 37244 34670 37256
rect 34900 37253 34928 37284
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 34664 37216 34897 37244
rect 34664 37204 34670 37216
rect 34885 37213 34897 37216
rect 34931 37213 34943 37247
rect 34885 37207 34943 37213
rect 34977 37247 35035 37253
rect 34977 37213 34989 37247
rect 35023 37244 35035 37247
rect 35986 37244 35992 37256
rect 35023 37216 35992 37244
rect 35023 37213 35035 37216
rect 34977 37207 35035 37213
rect 33778 37176 33784 37188
rect 33192 37148 33456 37176
rect 33739 37148 33784 37176
rect 33192 37136 33198 37148
rect 33778 37136 33784 37148
rect 33836 37136 33842 37188
rect 33870 37136 33876 37188
rect 33928 37176 33934 37188
rect 34992 37176 35020 37207
rect 35986 37204 35992 37216
rect 36044 37204 36050 37256
rect 36188 37253 36216 37284
rect 36722 37272 36728 37284
rect 36780 37272 36786 37324
rect 38197 37315 38255 37321
rect 38197 37281 38209 37315
rect 38243 37312 38255 37315
rect 38378 37312 38384 37324
rect 38243 37284 38384 37312
rect 38243 37281 38255 37284
rect 38197 37275 38255 37281
rect 38378 37272 38384 37284
rect 38436 37272 38442 37324
rect 38473 37315 38531 37321
rect 38473 37281 38485 37315
rect 38519 37312 38531 37315
rect 38519 37284 38976 37312
rect 38519 37281 38531 37284
rect 38473 37275 38531 37281
rect 36173 37247 36231 37253
rect 36173 37213 36185 37247
rect 36219 37213 36231 37247
rect 36354 37244 36360 37256
rect 36315 37216 36360 37244
rect 36173 37207 36231 37213
rect 36354 37204 36360 37216
rect 36412 37204 36418 37256
rect 36630 37244 36636 37256
rect 36591 37216 36636 37244
rect 36630 37204 36636 37216
rect 36688 37204 36694 37256
rect 37734 37204 37740 37256
rect 37792 37244 37798 37256
rect 38289 37247 38347 37253
rect 38289 37244 38301 37247
rect 37792 37216 38301 37244
rect 37792 37204 37798 37216
rect 38289 37213 38301 37216
rect 38335 37213 38347 37247
rect 38948 37244 38976 37284
rect 39022 37272 39028 37324
rect 39080 37312 39086 37324
rect 39080 37284 39125 37312
rect 39080 37272 39086 37284
rect 39574 37272 39580 37324
rect 39632 37312 39638 37324
rect 43346 37312 43352 37324
rect 39632 37284 40356 37312
rect 39632 37272 39638 37284
rect 39117 37247 39175 37253
rect 39117 37244 39129 37247
rect 38948 37216 39129 37244
rect 38289 37207 38347 37213
rect 39117 37213 39129 37216
rect 39163 37213 39175 37247
rect 40034 37244 40040 37256
rect 39995 37216 40040 37244
rect 39117 37207 39175 37213
rect 40034 37204 40040 37216
rect 40092 37204 40098 37256
rect 40328 37253 40356 37284
rect 42168 37284 42472 37312
rect 43307 37284 43352 37312
rect 40221 37247 40279 37253
rect 40221 37213 40233 37247
rect 40267 37213 40279 37247
rect 40221 37207 40279 37213
rect 40313 37247 40371 37253
rect 40313 37213 40325 37247
rect 40359 37213 40371 37247
rect 40313 37207 40371 37213
rect 40497 37247 40555 37253
rect 40497 37213 40509 37247
rect 40543 37244 40555 37247
rect 40586 37244 40592 37256
rect 40543 37216 40592 37244
rect 40543 37213 40555 37216
rect 40497 37207 40555 37213
rect 33928 37148 35020 37176
rect 35161 37179 35219 37185
rect 33928 37136 33934 37148
rect 35161 37145 35173 37179
rect 35207 37145 35219 37179
rect 35161 37139 35219 37145
rect 36817 37179 36875 37185
rect 36817 37145 36829 37179
rect 36863 37176 36875 37179
rect 39206 37176 39212 37188
rect 36863 37148 39212 37176
rect 36863 37145 36875 37148
rect 36817 37139 36875 37145
rect 34422 37108 34428 37120
rect 33060 37080 34428 37108
rect 29825 37071 29883 37077
rect 34422 37068 34428 37080
rect 34480 37108 34486 37120
rect 35176 37108 35204 37139
rect 39206 37136 39212 37148
rect 39264 37136 39270 37188
rect 39942 37136 39948 37188
rect 40000 37176 40006 37188
rect 40236 37176 40264 37207
rect 40586 37204 40592 37216
rect 40644 37204 40650 37256
rect 41506 37244 41512 37256
rect 41467 37216 41512 37244
rect 41506 37204 41512 37216
rect 41564 37204 41570 37256
rect 41782 37244 41788 37256
rect 41743 37216 41788 37244
rect 41782 37204 41788 37216
rect 41840 37244 41846 37256
rect 42168 37244 42196 37284
rect 41840 37216 42196 37244
rect 41840 37204 41846 37216
rect 42242 37204 42248 37256
rect 42300 37244 42306 37256
rect 42444 37253 42472 37284
rect 43346 37272 43352 37284
rect 43404 37272 43410 37324
rect 47504 37312 47532 37352
rect 47765 37349 47777 37383
rect 47811 37349 47823 37383
rect 47765 37343 47823 37349
rect 47504 37284 47624 37312
rect 42429 37247 42487 37253
rect 42300 37216 42345 37244
rect 42300 37204 42306 37216
rect 42429 37213 42441 37247
rect 42475 37213 42487 37247
rect 43438 37244 43444 37256
rect 43399 37216 43444 37244
rect 42429 37207 42487 37213
rect 43438 37204 43444 37216
rect 43496 37204 43502 37256
rect 46014 37244 46020 37256
rect 45975 37216 46020 37244
rect 46014 37204 46020 37216
rect 46072 37204 46078 37256
rect 46106 37204 46112 37256
rect 46164 37244 46170 37256
rect 46293 37247 46351 37253
rect 46293 37244 46305 37247
rect 46164 37216 46305 37244
rect 46164 37204 46170 37216
rect 46293 37213 46305 37216
rect 46339 37213 46351 37247
rect 46293 37207 46351 37213
rect 46566 37204 46572 37256
rect 46624 37244 46630 37256
rect 46661 37247 46719 37253
rect 46661 37244 46673 37247
rect 46624 37216 46673 37244
rect 46624 37204 46630 37216
rect 46661 37213 46673 37216
rect 46707 37213 46719 37247
rect 46661 37207 46719 37213
rect 46934 37204 46940 37256
rect 46992 37244 46998 37256
rect 47596 37253 47624 37284
rect 47489 37247 47547 37253
rect 47489 37244 47501 37247
rect 46992 37216 47501 37244
rect 46992 37204 46998 37216
rect 47489 37213 47501 37216
rect 47535 37213 47547 37247
rect 47489 37207 47547 37213
rect 47581 37247 47639 37253
rect 47581 37213 47593 37247
rect 47627 37213 47639 37247
rect 47780 37244 47808 37343
rect 49326 37340 49332 37392
rect 49384 37380 49390 37392
rect 51994 37380 52000 37392
rect 49384 37352 52000 37380
rect 49384 37340 49390 37352
rect 51994 37340 52000 37352
rect 52052 37340 52058 37392
rect 52914 37340 52920 37392
rect 52972 37380 52978 37392
rect 52972 37352 53420 37380
rect 52972 37340 52978 37352
rect 48590 37272 48596 37324
rect 48648 37272 48654 37324
rect 49421 37315 49479 37321
rect 49421 37281 49433 37315
rect 49467 37312 49479 37315
rect 50246 37312 50252 37324
rect 49467 37284 50252 37312
rect 49467 37281 49479 37284
rect 49421 37275 49479 37281
rect 50246 37272 50252 37284
rect 50304 37272 50310 37324
rect 51721 37315 51779 37321
rect 51721 37281 51733 37315
rect 51767 37312 51779 37315
rect 53282 37312 53288 37324
rect 51767 37284 53288 37312
rect 51767 37281 51779 37284
rect 51721 37275 51779 37281
rect 53282 37272 53288 37284
rect 53340 37272 53346 37324
rect 48225 37247 48283 37253
rect 48225 37244 48237 37247
rect 47780 37216 48237 37244
rect 47581 37207 47639 37213
rect 48225 37213 48237 37216
rect 48271 37213 48283 37247
rect 48225 37207 48283 37213
rect 40000 37148 40264 37176
rect 41693 37179 41751 37185
rect 40000 37136 40006 37148
rect 41693 37145 41705 37179
rect 41739 37176 41751 37179
rect 42702 37176 42708 37188
rect 41739 37148 42708 37176
rect 41739 37145 41751 37148
rect 41693 37139 41751 37145
rect 42702 37136 42708 37148
rect 42760 37136 42766 37188
rect 34480 37080 35204 37108
rect 34480 37068 34486 37080
rect 35618 37068 35624 37120
rect 35676 37108 35682 37120
rect 37458 37108 37464 37120
rect 35676 37080 37464 37108
rect 35676 37068 35682 37080
rect 37458 37068 37464 37080
rect 37516 37068 37522 37120
rect 37826 37108 37832 37120
rect 37787 37080 37832 37108
rect 37826 37068 37832 37080
rect 37884 37068 37890 37120
rect 40681 37111 40739 37117
rect 40681 37077 40693 37111
rect 40727 37108 40739 37111
rect 42518 37108 42524 37120
rect 40727 37080 42524 37108
rect 40727 37077 40739 37080
rect 40681 37071 40739 37077
rect 42518 37068 42524 37080
rect 42576 37068 42582 37120
rect 42613 37111 42671 37117
rect 42613 37077 42625 37111
rect 42659 37108 42671 37111
rect 45002 37108 45008 37120
rect 42659 37080 45008 37108
rect 42659 37077 42671 37080
rect 42613 37071 42671 37077
rect 45002 37068 45008 37080
rect 45060 37068 45066 37120
rect 45094 37068 45100 37120
rect 45152 37108 45158 37120
rect 45281 37111 45339 37117
rect 45281 37108 45293 37111
rect 45152 37080 45293 37108
rect 45152 37068 45158 37080
rect 45281 37077 45293 37080
rect 45327 37108 45339 37111
rect 45462 37108 45468 37120
rect 45327 37080 45468 37108
rect 45327 37077 45339 37080
rect 45281 37071 45339 37077
rect 45462 37068 45468 37080
rect 45520 37068 45526 37120
rect 47596 37108 47624 37207
rect 48314 37204 48320 37256
rect 48372 37244 48378 37256
rect 48608 37244 48636 37272
rect 48690 37247 48748 37253
rect 48690 37244 48702 37247
rect 48372 37216 48417 37244
rect 48608 37216 48702 37244
rect 48372 37204 48378 37216
rect 48690 37213 48702 37216
rect 48736 37213 48748 37247
rect 49326 37244 49332 37256
rect 49287 37216 49332 37244
rect 48690 37207 48748 37213
rect 49326 37204 49332 37216
rect 49384 37204 49390 37256
rect 49513 37247 49571 37253
rect 49513 37213 49525 37247
rect 49559 37213 49571 37247
rect 49513 37207 49571 37213
rect 47762 37176 47768 37188
rect 47723 37148 47768 37176
rect 47762 37136 47768 37148
rect 47820 37136 47826 37188
rect 48406 37136 48412 37188
rect 48464 37176 48470 37188
rect 48501 37179 48559 37185
rect 48501 37176 48513 37179
rect 48464 37148 48513 37176
rect 48464 37136 48470 37148
rect 48501 37145 48513 37148
rect 48547 37145 48559 37179
rect 48501 37139 48559 37145
rect 48593 37179 48651 37185
rect 48593 37145 48605 37179
rect 48639 37145 48651 37179
rect 49528 37176 49556 37207
rect 49694 37204 49700 37256
rect 49752 37244 49758 37256
rect 50709 37247 50767 37253
rect 50709 37244 50721 37247
rect 49752 37216 50721 37244
rect 49752 37204 49758 37216
rect 50709 37213 50721 37216
rect 50755 37213 50767 37247
rect 50709 37207 50767 37213
rect 50798 37204 50804 37256
rect 50856 37244 50862 37256
rect 50893 37247 50951 37253
rect 50893 37244 50905 37247
rect 50856 37216 50905 37244
rect 50856 37204 50862 37216
rect 50893 37213 50905 37216
rect 50939 37213 50951 37247
rect 50893 37207 50951 37213
rect 50982 37204 50988 37256
rect 51040 37244 51046 37256
rect 53392 37253 53420 37352
rect 54110 37340 54116 37392
rect 54168 37380 54174 37392
rect 54478 37380 54484 37392
rect 54168 37352 54484 37380
rect 54168 37340 54174 37352
rect 54478 37340 54484 37352
rect 54536 37340 54542 37392
rect 53558 37272 53564 37324
rect 53616 37312 53622 37324
rect 53653 37315 53711 37321
rect 53653 37312 53665 37315
rect 53616 37284 53665 37312
rect 53616 37272 53622 37284
rect 53653 37281 53665 37284
rect 53699 37281 53711 37315
rect 53653 37275 53711 37281
rect 54036 37284 54432 37312
rect 53377 37247 53435 37253
rect 51040 37238 53144 37244
rect 51040 37216 53328 37238
rect 51040 37204 51046 37216
rect 53116 37210 53328 37216
rect 50338 37176 50344 37188
rect 49528 37148 50344 37176
rect 48593 37139 48651 37145
rect 47854 37108 47860 37120
rect 47596 37080 47860 37108
rect 47854 37068 47860 37080
rect 47912 37108 47918 37120
rect 48608 37108 48636 37139
rect 50338 37136 50344 37148
rect 50396 37176 50402 37188
rect 52454 37176 52460 37188
rect 50396 37148 52460 37176
rect 50396 37136 50402 37148
rect 52454 37136 52460 37148
rect 52512 37136 52518 37188
rect 48682 37108 48688 37120
rect 47912 37080 48688 37108
rect 47912 37068 47918 37080
rect 48682 37068 48688 37080
rect 48740 37068 48746 37120
rect 48869 37111 48927 37117
rect 48869 37077 48881 37111
rect 48915 37108 48927 37111
rect 49142 37108 49148 37120
rect 48915 37080 49148 37108
rect 48915 37077 48927 37080
rect 48869 37071 48927 37077
rect 49142 37068 49148 37080
rect 49200 37068 49206 37120
rect 51994 37068 52000 37120
rect 52052 37108 52058 37120
rect 52273 37111 52331 37117
rect 52273 37108 52285 37111
rect 52052 37080 52285 37108
rect 52052 37068 52058 37080
rect 52273 37077 52285 37080
rect 52319 37108 52331 37111
rect 52733 37111 52791 37117
rect 52733 37108 52745 37111
rect 52319 37080 52745 37108
rect 52319 37077 52331 37080
rect 52273 37071 52331 37077
rect 52733 37077 52745 37080
rect 52779 37108 52791 37111
rect 53190 37108 53196 37120
rect 52779 37080 53196 37108
rect 52779 37077 52791 37080
rect 52733 37071 52791 37077
rect 53190 37068 53196 37080
rect 53248 37068 53254 37120
rect 53300 37108 53328 37210
rect 53377 37213 53389 37247
rect 53423 37244 53435 37247
rect 54036 37244 54064 37284
rect 53423 37216 54064 37244
rect 54113 37247 54171 37253
rect 53423 37213 53435 37216
rect 53377 37207 53435 37213
rect 54113 37213 54125 37247
rect 54159 37213 54171 37247
rect 54113 37207 54171 37213
rect 53653 37179 53711 37185
rect 53653 37145 53665 37179
rect 53699 37176 53711 37179
rect 54128 37176 54156 37207
rect 54202 37204 54208 37256
rect 54260 37244 54266 37256
rect 54404 37244 54432 37284
rect 55858 37272 55864 37324
rect 55916 37312 55922 37324
rect 55953 37315 56011 37321
rect 55953 37312 55965 37315
rect 55916 37284 55965 37312
rect 55916 37272 55922 37284
rect 55953 37281 55965 37284
rect 55999 37281 56011 37315
rect 55953 37275 56011 37281
rect 54481 37247 54539 37253
rect 54481 37244 54493 37247
rect 54260 37216 54305 37244
rect 54404 37216 54493 37244
rect 54260 37204 54266 37216
rect 54481 37213 54493 37216
rect 54527 37213 54539 37247
rect 54481 37207 54539 37213
rect 54570 37204 54576 37256
rect 54628 37253 54634 37256
rect 54628 37244 54636 37253
rect 54628 37216 54673 37244
rect 54628 37207 54636 37216
rect 54628 37204 54634 37207
rect 55766 37204 55772 37256
rect 55824 37244 55830 37256
rect 56045 37247 56103 37253
rect 56045 37244 56057 37247
rect 55824 37216 56057 37244
rect 55824 37204 55830 37216
rect 56045 37213 56057 37216
rect 56091 37213 56103 37247
rect 56045 37207 56103 37213
rect 54386 37176 54392 37188
rect 53699 37148 54156 37176
rect 54299 37148 54392 37176
rect 53699 37145 53711 37148
rect 53653 37139 53711 37145
rect 54386 37136 54392 37148
rect 54444 37136 54450 37188
rect 54404 37108 54432 37136
rect 53300 37080 54432 37108
rect 54757 37111 54815 37117
rect 54757 37077 54769 37111
rect 54803 37108 54815 37111
rect 54846 37108 54852 37120
rect 54803 37080 54852 37108
rect 54803 37077 54815 37080
rect 54757 37071 54815 37077
rect 54846 37068 54852 37080
rect 54904 37068 54910 37120
rect 57974 37108 57980 37120
rect 57935 37080 57980 37108
rect 57974 37068 57980 37080
rect 58032 37068 58038 37120
rect 1104 37018 58880 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 58880 37018
rect 1104 36944 58880 36966
rect 28258 36864 28264 36916
rect 28316 36904 28322 36916
rect 29730 36904 29736 36916
rect 28316 36876 29736 36904
rect 28316 36864 28322 36876
rect 29730 36864 29736 36876
rect 29788 36864 29794 36916
rect 30006 36904 30012 36916
rect 29967 36876 30012 36904
rect 30006 36864 30012 36876
rect 30064 36864 30070 36916
rect 33778 36864 33784 36916
rect 33836 36904 33842 36916
rect 34333 36907 34391 36913
rect 34333 36904 34345 36907
rect 33836 36876 34345 36904
rect 33836 36864 33842 36876
rect 34333 36873 34345 36876
rect 34379 36904 34391 36907
rect 35802 36904 35808 36916
rect 34379 36876 35808 36904
rect 34379 36873 34391 36876
rect 34333 36867 34391 36873
rect 35802 36864 35808 36876
rect 35860 36864 35866 36916
rect 35989 36907 36047 36913
rect 35989 36873 36001 36907
rect 36035 36904 36047 36907
rect 36630 36904 36636 36916
rect 36035 36876 36636 36904
rect 36035 36873 36047 36876
rect 35989 36867 36047 36873
rect 36630 36864 36636 36876
rect 36688 36864 36694 36916
rect 38473 36907 38531 36913
rect 38473 36873 38485 36907
rect 38519 36904 38531 36907
rect 39022 36904 39028 36916
rect 38519 36876 39028 36904
rect 38519 36873 38531 36876
rect 38473 36867 38531 36873
rect 39022 36864 39028 36876
rect 39080 36864 39086 36916
rect 39206 36864 39212 36916
rect 39264 36904 39270 36916
rect 43530 36904 43536 36916
rect 39264 36876 43536 36904
rect 39264 36864 39270 36876
rect 43530 36864 43536 36876
rect 43588 36864 43594 36916
rect 48225 36907 48283 36913
rect 45572 36876 48176 36904
rect 28997 36839 29055 36845
rect 28997 36805 29009 36839
rect 29043 36836 29055 36839
rect 30190 36836 30196 36848
rect 29043 36808 30196 36836
rect 29043 36805 29055 36808
rect 28997 36799 29055 36805
rect 30190 36796 30196 36808
rect 30248 36796 30254 36848
rect 31386 36836 31392 36848
rect 30484 36808 31392 36836
rect 28166 36728 28172 36780
rect 28224 36768 28230 36780
rect 28902 36768 28908 36780
rect 28224 36740 28908 36768
rect 28224 36728 28230 36740
rect 28902 36728 28908 36740
rect 28960 36728 28966 36780
rect 29086 36728 29092 36780
rect 29144 36768 29150 36780
rect 29181 36771 29239 36777
rect 29181 36768 29193 36771
rect 29144 36740 29193 36768
rect 29144 36728 29150 36740
rect 29181 36737 29193 36740
rect 29227 36737 29239 36771
rect 29914 36768 29920 36780
rect 29875 36740 29920 36768
rect 29181 36731 29239 36737
rect 29914 36728 29920 36740
rect 29972 36728 29978 36780
rect 30484 36768 30512 36808
rect 30208 36740 30512 36768
rect 29362 36660 29368 36712
rect 29420 36700 29426 36712
rect 30208 36700 30236 36740
rect 30558 36728 30564 36780
rect 30616 36768 30622 36780
rect 30745 36771 30803 36777
rect 30745 36768 30757 36771
rect 30616 36740 30757 36768
rect 30616 36728 30622 36740
rect 30745 36737 30757 36740
rect 30791 36737 30803 36771
rect 30745 36731 30803 36737
rect 30926 36728 30932 36780
rect 30984 36768 30990 36780
rect 31220 36777 31248 36808
rect 31386 36796 31392 36808
rect 31444 36796 31450 36848
rect 32493 36839 32551 36845
rect 32493 36805 32505 36839
rect 32539 36836 32551 36839
rect 32858 36836 32864 36848
rect 32539 36808 32864 36836
rect 32539 36805 32551 36808
rect 32493 36799 32551 36805
rect 32858 36796 32864 36808
rect 32916 36796 32922 36848
rect 32950 36796 32956 36848
rect 33008 36836 33014 36848
rect 37826 36836 37832 36848
rect 33008 36808 34652 36836
rect 33008 36796 33014 36808
rect 34624 36780 34652 36808
rect 35452 36808 37832 36836
rect 31113 36771 31171 36777
rect 31113 36768 31125 36771
rect 30984 36740 31125 36768
rect 30984 36728 30990 36740
rect 31113 36737 31125 36740
rect 31159 36737 31171 36771
rect 31113 36731 31171 36737
rect 31205 36771 31263 36777
rect 31205 36737 31217 36771
rect 31251 36737 31263 36771
rect 32674 36768 32680 36780
rect 32635 36740 32680 36768
rect 31205 36731 31263 36737
rect 32674 36728 32680 36740
rect 32732 36728 32738 36780
rect 32766 36728 32772 36780
rect 32824 36768 32830 36780
rect 33321 36771 33379 36777
rect 33321 36768 33333 36771
rect 32824 36740 33333 36768
rect 32824 36728 32830 36740
rect 33321 36737 33333 36740
rect 33367 36737 33379 36771
rect 34422 36768 34428 36780
rect 34335 36740 34428 36768
rect 33321 36731 33379 36737
rect 34422 36728 34428 36740
rect 34480 36728 34486 36780
rect 34606 36728 34612 36780
rect 34664 36768 34670 36780
rect 35345 36771 35403 36777
rect 35345 36768 35357 36771
rect 34664 36740 35357 36768
rect 34664 36728 34670 36740
rect 35345 36737 35357 36740
rect 35391 36737 35403 36771
rect 35345 36731 35403 36737
rect 29420 36672 30236 36700
rect 29420 36660 29426 36672
rect 30374 36660 30380 36712
rect 30432 36700 30438 36712
rect 30650 36700 30656 36712
rect 30432 36672 30656 36700
rect 30432 36660 30438 36672
rect 30650 36660 30656 36672
rect 30708 36660 30714 36712
rect 34238 36700 34244 36712
rect 34199 36672 34244 36700
rect 34238 36660 34244 36672
rect 34296 36660 34302 36712
rect 29178 36632 29184 36644
rect 29139 36604 29184 36632
rect 29178 36592 29184 36604
rect 29236 36592 29242 36644
rect 29270 36592 29276 36644
rect 29328 36632 29334 36644
rect 29328 36604 33548 36632
rect 29328 36592 29334 36604
rect 32861 36567 32919 36573
rect 32861 36533 32873 36567
rect 32907 36564 32919 36567
rect 33134 36564 33140 36576
rect 32907 36536 33140 36564
rect 32907 36533 32919 36536
rect 32861 36527 32919 36533
rect 33134 36524 33140 36536
rect 33192 36524 33198 36576
rect 33520 36573 33548 36604
rect 33505 36567 33563 36573
rect 33505 36533 33517 36567
rect 33551 36564 33563 36567
rect 33962 36564 33968 36576
rect 33551 36536 33968 36564
rect 33551 36533 33563 36536
rect 33505 36527 33563 36533
rect 33962 36524 33968 36536
rect 34020 36524 34026 36576
rect 34440 36564 34468 36728
rect 34793 36635 34851 36641
rect 34793 36601 34805 36635
rect 34839 36632 34851 36635
rect 35452 36632 35480 36808
rect 37826 36796 37832 36808
rect 37884 36796 37890 36848
rect 40034 36836 40040 36848
rect 39040 36808 40040 36836
rect 35529 36771 35587 36777
rect 35529 36737 35541 36771
rect 35575 36737 35587 36771
rect 35529 36731 35587 36737
rect 35621 36771 35679 36777
rect 35621 36737 35633 36771
rect 35667 36737 35679 36771
rect 35621 36731 35679 36737
rect 35713 36771 35771 36777
rect 35713 36737 35725 36771
rect 35759 36768 35771 36771
rect 35986 36768 35992 36780
rect 35759 36740 35992 36768
rect 35759 36737 35771 36740
rect 35713 36731 35771 36737
rect 34839 36604 35480 36632
rect 34839 36601 34851 36604
rect 34793 36595 34851 36601
rect 35544 36564 35572 36731
rect 35636 36632 35664 36731
rect 35986 36728 35992 36740
rect 36044 36768 36050 36780
rect 36449 36771 36507 36777
rect 36449 36768 36461 36771
rect 36044 36740 36461 36768
rect 36044 36728 36050 36740
rect 36449 36737 36461 36740
rect 36495 36737 36507 36771
rect 36449 36731 36507 36737
rect 36633 36771 36691 36777
rect 36633 36737 36645 36771
rect 36679 36768 36691 36771
rect 37182 36768 37188 36780
rect 36679 36740 37188 36768
rect 36679 36737 36691 36740
rect 36633 36731 36691 36737
rect 35802 36660 35808 36712
rect 35860 36700 35866 36712
rect 36541 36703 36599 36709
rect 36541 36700 36553 36703
rect 35860 36672 36553 36700
rect 35860 36660 35866 36672
rect 36541 36669 36553 36672
rect 36587 36669 36599 36703
rect 36541 36663 36599 36669
rect 36170 36632 36176 36644
rect 35636 36604 36176 36632
rect 36170 36592 36176 36604
rect 36228 36592 36234 36644
rect 36648 36564 36676 36731
rect 37182 36728 37188 36740
rect 37240 36728 37246 36780
rect 38102 36768 38108 36780
rect 38063 36740 38108 36768
rect 38102 36728 38108 36740
rect 38160 36728 38166 36780
rect 38930 36768 38936 36780
rect 38891 36740 38936 36768
rect 38930 36728 38936 36740
rect 38988 36728 38994 36780
rect 39040 36777 39068 36808
rect 40034 36796 40040 36808
rect 40092 36836 40098 36848
rect 44082 36836 44088 36848
rect 40092 36808 41184 36836
rect 40092 36796 40098 36808
rect 39025 36771 39083 36777
rect 39025 36737 39037 36771
rect 39071 36737 39083 36771
rect 39025 36731 39083 36737
rect 39117 36771 39175 36777
rect 39117 36737 39129 36771
rect 39163 36737 39175 36771
rect 39117 36731 39175 36737
rect 38010 36700 38016 36712
rect 37971 36672 38016 36700
rect 38010 36660 38016 36672
rect 38068 36660 38074 36712
rect 39132 36700 39160 36731
rect 39206 36728 39212 36780
rect 39264 36768 39270 36780
rect 39577 36771 39635 36777
rect 39577 36768 39589 36771
rect 39264 36740 39589 36768
rect 39264 36728 39270 36740
rect 39577 36737 39589 36740
rect 39623 36768 39635 36771
rect 39942 36768 39948 36780
rect 39623 36740 39948 36768
rect 39623 36737 39635 36740
rect 39577 36731 39635 36737
rect 39942 36728 39948 36740
rect 40000 36728 40006 36780
rect 40218 36768 40224 36780
rect 40179 36740 40224 36768
rect 40218 36728 40224 36740
rect 40276 36728 40282 36780
rect 41156 36777 41184 36808
rect 41616 36808 44088 36836
rect 41141 36771 41199 36777
rect 41141 36737 41153 36771
rect 41187 36737 41199 36771
rect 41414 36768 41420 36780
rect 41375 36740 41420 36768
rect 41141 36731 41199 36737
rect 41414 36728 41420 36740
rect 41472 36728 41478 36780
rect 41616 36777 41644 36808
rect 44082 36796 44088 36808
rect 44140 36796 44146 36848
rect 41601 36771 41659 36777
rect 41601 36737 41613 36771
rect 41647 36737 41659 36771
rect 42886 36768 42892 36780
rect 42847 36740 42892 36768
rect 41601 36731 41659 36737
rect 42886 36728 42892 36740
rect 42944 36728 42950 36780
rect 44266 36728 44272 36780
rect 44324 36768 44330 36780
rect 44637 36771 44695 36777
rect 44637 36768 44649 36771
rect 44324 36740 44649 36768
rect 44324 36728 44330 36740
rect 44637 36737 44649 36740
rect 44683 36737 44695 36771
rect 44637 36731 44695 36737
rect 45186 36728 45192 36780
rect 45244 36768 45250 36780
rect 45281 36771 45339 36777
rect 45281 36768 45293 36771
rect 45244 36740 45293 36768
rect 45244 36728 45250 36740
rect 45281 36737 45293 36740
rect 45327 36737 45339 36771
rect 45462 36768 45468 36780
rect 45423 36740 45468 36768
rect 45281 36731 45339 36737
rect 45462 36728 45468 36740
rect 45520 36728 45526 36780
rect 45572 36777 45600 36876
rect 46661 36839 46719 36845
rect 46661 36805 46673 36839
rect 46707 36836 46719 36839
rect 47762 36836 47768 36848
rect 46707 36808 47768 36836
rect 46707 36805 46719 36808
rect 46661 36799 46719 36805
rect 47762 36796 47768 36808
rect 47820 36796 47826 36848
rect 48148 36836 48176 36876
rect 48225 36873 48237 36907
rect 48271 36904 48283 36907
rect 48590 36904 48596 36916
rect 48271 36876 48596 36904
rect 48271 36873 48283 36876
rect 48225 36867 48283 36873
rect 48590 36864 48596 36876
rect 48648 36864 48654 36916
rect 50062 36864 50068 36916
rect 50120 36904 50126 36916
rect 50157 36907 50215 36913
rect 50157 36904 50169 36907
rect 50120 36876 50169 36904
rect 50120 36864 50126 36876
rect 50157 36873 50169 36876
rect 50203 36904 50215 36907
rect 50706 36904 50712 36916
rect 50203 36876 50712 36904
rect 50203 36873 50215 36876
rect 50157 36867 50215 36873
rect 50706 36864 50712 36876
rect 50764 36864 50770 36916
rect 51445 36907 51503 36913
rect 51445 36873 51457 36907
rect 51491 36904 51503 36907
rect 52362 36904 52368 36916
rect 51491 36876 52368 36904
rect 51491 36873 51503 36876
rect 51445 36867 51503 36873
rect 49970 36836 49976 36848
rect 48148 36808 49976 36836
rect 49970 36796 49976 36808
rect 50028 36796 50034 36848
rect 50338 36836 50344 36848
rect 50299 36808 50344 36836
rect 50338 36796 50344 36808
rect 50396 36796 50402 36848
rect 51920 36845 51948 36876
rect 52362 36864 52368 36876
rect 52420 36904 52426 36916
rect 52914 36904 52920 36916
rect 52420 36876 52920 36904
rect 52420 36864 52426 36876
rect 52914 36864 52920 36876
rect 52972 36904 52978 36916
rect 56137 36907 56195 36913
rect 56137 36904 56149 36907
rect 52972 36876 56149 36904
rect 52972 36864 52978 36876
rect 56137 36873 56149 36876
rect 56183 36873 56195 36907
rect 56137 36867 56195 36873
rect 51905 36839 51963 36845
rect 51905 36805 51917 36839
rect 51951 36805 51963 36839
rect 51905 36799 51963 36805
rect 51994 36796 52000 36848
rect 52052 36836 52058 36848
rect 52181 36839 52239 36845
rect 52181 36836 52193 36839
rect 52052 36808 52193 36836
rect 52052 36796 52058 36808
rect 52181 36805 52193 36808
rect 52227 36805 52239 36839
rect 53466 36836 53472 36848
rect 52181 36799 52239 36805
rect 53300 36808 53472 36836
rect 45557 36771 45615 36777
rect 45557 36737 45569 36771
rect 45603 36737 45615 36771
rect 45557 36731 45615 36737
rect 46014 36728 46020 36780
rect 46072 36768 46078 36780
rect 46290 36768 46296 36780
rect 46072 36740 46296 36768
rect 46072 36728 46078 36740
rect 46290 36728 46296 36740
rect 46348 36768 46354 36780
rect 46385 36771 46443 36777
rect 46385 36768 46397 36771
rect 46348 36740 46397 36768
rect 46348 36728 46354 36740
rect 46385 36737 46397 36740
rect 46431 36737 46443 36771
rect 46385 36731 46443 36737
rect 46566 36728 46572 36780
rect 46624 36768 46630 36780
rect 46753 36771 46811 36777
rect 46753 36768 46765 36771
rect 46624 36740 46765 36768
rect 46624 36728 46630 36740
rect 46753 36737 46765 36740
rect 46799 36737 46811 36771
rect 49234 36768 49240 36780
rect 49195 36740 49240 36768
rect 46753 36731 46811 36737
rect 49234 36728 49240 36740
rect 49292 36728 49298 36780
rect 50065 36771 50123 36777
rect 50065 36737 50077 36771
rect 50111 36737 50123 36771
rect 52086 36768 52092 36780
rect 52047 36740 52092 36768
rect 50065 36731 50123 36737
rect 39040 36672 39160 36700
rect 36722 36592 36728 36644
rect 36780 36632 36786 36644
rect 39040 36632 39068 36672
rect 42978 36660 42984 36712
rect 43036 36700 43042 36712
rect 43036 36672 43116 36700
rect 43036 36660 43042 36672
rect 39482 36632 39488 36644
rect 36780 36604 39488 36632
rect 36780 36592 36786 36604
rect 39482 36592 39488 36604
rect 39540 36632 39546 36644
rect 40405 36635 40463 36641
rect 40405 36632 40417 36635
rect 39540 36604 40417 36632
rect 39540 36592 39546 36604
rect 40405 36601 40417 36604
rect 40451 36601 40463 36635
rect 40405 36595 40463 36601
rect 34440 36536 36676 36564
rect 38010 36524 38016 36576
rect 38068 36564 38074 36576
rect 38378 36564 38384 36576
rect 38068 36536 38384 36564
rect 38068 36524 38074 36536
rect 38378 36524 38384 36536
rect 38436 36524 38442 36576
rect 39206 36524 39212 36576
rect 39264 36564 39270 36576
rect 39669 36567 39727 36573
rect 39669 36564 39681 36567
rect 39264 36536 39681 36564
rect 39264 36524 39270 36536
rect 39669 36533 39681 36536
rect 39715 36564 39727 36567
rect 40586 36564 40592 36576
rect 39715 36536 40592 36564
rect 39715 36533 39727 36536
rect 39669 36527 39727 36533
rect 40586 36524 40592 36536
rect 40644 36524 40650 36576
rect 40957 36567 41015 36573
rect 40957 36533 40969 36567
rect 41003 36564 41015 36567
rect 42978 36564 42984 36576
rect 41003 36536 42984 36564
rect 41003 36533 41015 36536
rect 40957 36527 41015 36533
rect 42978 36524 42984 36536
rect 43036 36524 43042 36576
rect 43088 36573 43116 36672
rect 44174 36660 44180 36712
rect 44232 36700 44238 36712
rect 44453 36703 44511 36709
rect 44453 36700 44465 36703
rect 44232 36672 44465 36700
rect 44232 36660 44238 36672
rect 44453 36669 44465 36672
rect 44499 36700 44511 36703
rect 46106 36700 46112 36712
rect 44499 36672 46112 36700
rect 44499 36669 44511 36672
rect 44453 36663 44511 36669
rect 46106 36660 46112 36672
rect 46164 36700 46170 36712
rect 46201 36703 46259 36709
rect 46201 36700 46213 36703
rect 46164 36672 46213 36700
rect 46164 36660 46170 36672
rect 46201 36669 46213 36672
rect 46247 36669 46259 36703
rect 46842 36700 46848 36712
rect 46201 36663 46259 36669
rect 46308 36672 46848 36700
rect 44821 36635 44879 36641
rect 44821 36601 44833 36635
rect 44867 36632 44879 36635
rect 46308 36632 46336 36672
rect 46842 36660 46848 36672
rect 46900 36700 46906 36712
rect 47765 36703 47823 36709
rect 47765 36700 47777 36703
rect 46900 36672 47777 36700
rect 46900 36660 46906 36672
rect 47765 36669 47777 36672
rect 47811 36669 47823 36703
rect 49142 36700 49148 36712
rect 49103 36672 49148 36700
rect 47765 36663 47823 36669
rect 49142 36660 49148 36672
rect 49200 36660 49206 36712
rect 49605 36703 49663 36709
rect 49605 36669 49617 36703
rect 49651 36700 49663 36703
rect 49694 36700 49700 36712
rect 49651 36672 49700 36700
rect 49651 36669 49663 36672
rect 49605 36663 49663 36669
rect 49694 36660 49700 36672
rect 49752 36660 49758 36712
rect 48130 36632 48136 36644
rect 44867 36604 46336 36632
rect 48091 36604 48136 36632
rect 44867 36601 44879 36604
rect 44821 36595 44879 36601
rect 48130 36592 48136 36604
rect 48188 36592 48194 36644
rect 50080 36632 50108 36731
rect 52086 36728 52092 36740
rect 52144 36728 52150 36780
rect 52270 36768 52276 36780
rect 52328 36777 52334 36780
rect 52236 36740 52276 36768
rect 52270 36728 52276 36740
rect 52328 36731 52336 36777
rect 53190 36768 53196 36780
rect 53151 36740 53196 36768
rect 52328 36728 52334 36731
rect 53190 36728 53196 36740
rect 53248 36728 53254 36780
rect 53300 36777 53328 36808
rect 53466 36796 53472 36808
rect 53524 36796 53530 36848
rect 53285 36771 53343 36777
rect 53285 36737 53297 36771
rect 53331 36737 53343 36771
rect 53285 36731 53343 36737
rect 53377 36771 53435 36777
rect 53377 36737 53389 36771
rect 53423 36737 53435 36771
rect 53558 36768 53564 36780
rect 53471 36740 53564 36768
rect 53377 36731 53435 36737
rect 52181 36703 52239 36709
rect 52181 36669 52193 36703
rect 52227 36700 52239 36703
rect 53392 36700 53420 36731
rect 53558 36728 53564 36740
rect 53616 36728 53622 36780
rect 53650 36728 53656 36780
rect 53708 36768 53714 36780
rect 54757 36771 54815 36777
rect 54757 36768 54769 36771
rect 53708 36740 54769 36768
rect 53708 36728 53714 36740
rect 54757 36737 54769 36740
rect 54803 36737 54815 36771
rect 54757 36731 54815 36737
rect 52227 36672 53420 36700
rect 52227 36669 52239 36672
rect 52181 36663 52239 36669
rect 53576 36632 53604 36728
rect 54846 36700 54852 36712
rect 54807 36672 54852 36700
rect 54846 36660 54852 36672
rect 54904 36660 54910 36712
rect 50080 36604 53604 36632
rect 55677 36635 55735 36641
rect 55677 36601 55689 36635
rect 55723 36632 55735 36635
rect 56226 36632 56232 36644
rect 55723 36604 56232 36632
rect 55723 36601 55735 36604
rect 55677 36595 55735 36601
rect 56226 36592 56232 36604
rect 56284 36592 56290 36644
rect 43073 36567 43131 36573
rect 43073 36533 43085 36567
rect 43119 36564 43131 36567
rect 43990 36564 43996 36576
rect 43119 36536 43996 36564
rect 43119 36533 43131 36536
rect 43073 36527 43131 36533
rect 43990 36524 43996 36536
rect 44048 36524 44054 36576
rect 45094 36524 45100 36576
rect 45152 36564 45158 36576
rect 45281 36567 45339 36573
rect 45281 36564 45293 36567
rect 45152 36536 45293 36564
rect 45152 36524 45158 36536
rect 45281 36533 45293 36536
rect 45327 36533 45339 36567
rect 45281 36527 45339 36533
rect 46290 36524 46296 36576
rect 46348 36564 46354 36576
rect 47394 36564 47400 36576
rect 46348 36536 47400 36564
rect 46348 36524 46354 36536
rect 47394 36524 47400 36536
rect 47452 36524 47458 36576
rect 47578 36524 47584 36576
rect 47636 36564 47642 36576
rect 50062 36564 50068 36576
rect 47636 36536 50068 36564
rect 47636 36524 47642 36536
rect 50062 36524 50068 36536
rect 50120 36524 50126 36576
rect 50338 36564 50344 36576
rect 50299 36536 50344 36564
rect 50338 36524 50344 36536
rect 50396 36524 50402 36576
rect 50706 36524 50712 36576
rect 50764 36564 50770 36576
rect 50801 36567 50859 36573
rect 50801 36564 50813 36567
rect 50764 36536 50813 36564
rect 50764 36524 50770 36536
rect 50801 36533 50813 36536
rect 50847 36533 50859 36567
rect 50801 36527 50859 36533
rect 52822 36524 52828 36576
rect 52880 36564 52886 36576
rect 52917 36567 52975 36573
rect 52917 36564 52929 36567
rect 52880 36536 52929 36564
rect 52880 36524 52886 36536
rect 52917 36533 52929 36536
rect 52963 36533 52975 36567
rect 52917 36527 52975 36533
rect 54113 36567 54171 36573
rect 54113 36533 54125 36567
rect 54159 36564 54171 36567
rect 54202 36564 54208 36576
rect 54159 36536 54208 36564
rect 54159 36533 54171 36536
rect 54113 36527 54171 36533
rect 54202 36524 54208 36536
rect 54260 36564 54266 36576
rect 54754 36564 54760 36576
rect 54260 36536 54760 36564
rect 54260 36524 54266 36536
rect 54754 36524 54760 36536
rect 54812 36524 54818 36576
rect 55122 36564 55128 36576
rect 55083 36536 55128 36564
rect 55122 36524 55128 36536
rect 55180 36524 55186 36576
rect 56594 36524 56600 36576
rect 56652 36564 56658 36576
rect 56689 36567 56747 36573
rect 56689 36564 56701 36567
rect 56652 36536 56701 36564
rect 56652 36524 56658 36536
rect 56689 36533 56701 36536
rect 56735 36564 56747 36567
rect 57333 36567 57391 36573
rect 57333 36564 57345 36567
rect 56735 36536 57345 36564
rect 56735 36533 56747 36536
rect 56689 36527 56747 36533
rect 57333 36533 57345 36536
rect 57379 36564 57391 36567
rect 57974 36564 57980 36576
rect 57379 36536 57980 36564
rect 57379 36533 57391 36536
rect 57333 36527 57391 36533
rect 57974 36524 57980 36536
rect 58032 36564 58038 36576
rect 58069 36567 58127 36573
rect 58069 36564 58081 36567
rect 58032 36536 58081 36564
rect 58032 36524 58038 36536
rect 58069 36533 58081 36536
rect 58115 36533 58127 36567
rect 58069 36527 58127 36533
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 29181 36363 29239 36369
rect 29181 36329 29193 36363
rect 29227 36360 29239 36363
rect 29914 36360 29920 36372
rect 29227 36332 29920 36360
rect 29227 36329 29239 36332
rect 29181 36323 29239 36329
rect 29914 36320 29920 36332
rect 29972 36320 29978 36372
rect 33134 36320 33140 36372
rect 33192 36360 33198 36372
rect 34054 36360 34060 36372
rect 33192 36332 34060 36360
rect 33192 36320 33198 36332
rect 34054 36320 34060 36332
rect 34112 36320 34118 36372
rect 34238 36320 34244 36372
rect 34296 36360 34302 36372
rect 34885 36363 34943 36369
rect 34885 36360 34897 36363
rect 34296 36332 34897 36360
rect 34296 36320 34302 36332
rect 34885 36329 34897 36332
rect 34931 36329 34943 36363
rect 34885 36323 34943 36329
rect 36630 36320 36636 36372
rect 36688 36360 36694 36372
rect 40218 36360 40224 36372
rect 36688 36332 40224 36360
rect 36688 36320 36694 36332
rect 40218 36320 40224 36332
rect 40276 36320 40282 36372
rect 41233 36363 41291 36369
rect 41233 36329 41245 36363
rect 41279 36360 41291 36363
rect 41506 36360 41512 36372
rect 41279 36332 41512 36360
rect 41279 36329 41291 36332
rect 41233 36323 41291 36329
rect 41506 36320 41512 36332
rect 41564 36320 41570 36372
rect 44637 36363 44695 36369
rect 44637 36329 44649 36363
rect 44683 36360 44695 36363
rect 49234 36360 49240 36372
rect 44683 36332 49240 36360
rect 44683 36329 44695 36332
rect 44637 36323 44695 36329
rect 49234 36320 49240 36332
rect 49292 36320 49298 36372
rect 29822 36292 29828 36304
rect 29783 36264 29828 36292
rect 29822 36252 29828 36264
rect 29880 36252 29886 36304
rect 31478 36252 31484 36304
rect 31536 36292 31542 36304
rect 33686 36292 33692 36304
rect 31536 36264 33692 36292
rect 31536 36252 31542 36264
rect 33686 36252 33692 36264
rect 33744 36252 33750 36304
rect 33985 36264 38153 36292
rect 30374 36184 30380 36236
rect 30432 36224 30438 36236
rect 30469 36227 30527 36233
rect 30469 36224 30481 36227
rect 30432 36196 30481 36224
rect 30432 36184 30438 36196
rect 30469 36193 30481 36196
rect 30515 36193 30527 36227
rect 30926 36224 30932 36236
rect 30887 36196 30932 36224
rect 30469 36187 30527 36193
rect 30926 36184 30932 36196
rect 30984 36224 30990 36236
rect 31386 36224 31392 36236
rect 30984 36196 31392 36224
rect 30984 36184 30990 36196
rect 31386 36184 31392 36196
rect 31444 36224 31450 36236
rect 32861 36227 32919 36233
rect 31444 36196 31754 36224
rect 31444 36184 31450 36196
rect 28902 36156 28908 36168
rect 28863 36128 28908 36156
rect 28902 36116 28908 36128
rect 28960 36116 28966 36168
rect 29270 36116 29276 36168
rect 29328 36156 29334 36168
rect 29733 36159 29791 36165
rect 29733 36156 29745 36159
rect 29328 36128 29745 36156
rect 29328 36116 29334 36128
rect 29733 36125 29745 36128
rect 29779 36125 29791 36159
rect 30558 36156 30564 36168
rect 30519 36128 30564 36156
rect 29733 36119 29791 36125
rect 30558 36116 30564 36128
rect 30616 36116 30622 36168
rect 31021 36159 31079 36165
rect 31021 36125 31033 36159
rect 31067 36125 31079 36159
rect 31726 36156 31754 36196
rect 32861 36193 32873 36227
rect 32907 36224 32919 36227
rect 33042 36224 33048 36236
rect 32907 36196 33048 36224
rect 32907 36193 32919 36196
rect 32861 36187 32919 36193
rect 33042 36184 33048 36196
rect 33100 36224 33106 36236
rect 33985 36224 34013 36264
rect 33100 36196 34013 36224
rect 33100 36184 33106 36196
rect 32033 36159 32091 36165
rect 32033 36156 32045 36159
rect 31726 36128 32045 36156
rect 31021 36119 31079 36125
rect 32033 36125 32045 36128
rect 32079 36125 32091 36159
rect 33502 36156 33508 36168
rect 33463 36128 33508 36156
rect 32033 36119 32091 36125
rect 29178 36088 29184 36100
rect 29139 36060 29184 36088
rect 29178 36048 29184 36060
rect 29236 36048 29242 36100
rect 29822 36048 29828 36100
rect 29880 36088 29886 36100
rect 31036 36088 31064 36119
rect 33502 36116 33508 36128
rect 33560 36116 33566 36168
rect 33985 36165 34013 36196
rect 34054 36184 34060 36236
rect 34112 36224 34118 36236
rect 36081 36227 36139 36233
rect 36081 36224 36093 36227
rect 34112 36196 36093 36224
rect 34112 36184 34118 36196
rect 36081 36193 36093 36196
rect 36127 36193 36139 36227
rect 36722 36224 36728 36236
rect 36081 36187 36139 36193
rect 36556 36196 36728 36224
rect 33598 36159 33656 36165
rect 33598 36125 33610 36159
rect 33644 36125 33656 36159
rect 33598 36119 33656 36125
rect 33970 36159 34028 36165
rect 33970 36125 33982 36159
rect 34016 36125 34028 36159
rect 33970 36119 34028 36125
rect 35069 36159 35127 36165
rect 35069 36125 35081 36159
rect 35115 36125 35127 36159
rect 35069 36119 35127 36125
rect 35345 36159 35403 36165
rect 35345 36125 35357 36159
rect 35391 36156 35403 36159
rect 35986 36156 35992 36168
rect 35391 36128 35992 36156
rect 35391 36125 35403 36128
rect 35345 36119 35403 36125
rect 29880 36060 31064 36088
rect 29880 36048 29886 36060
rect 33318 36048 33324 36100
rect 33376 36088 33382 36100
rect 33612 36088 33640 36119
rect 33778 36088 33784 36100
rect 33376 36060 33640 36088
rect 33739 36060 33784 36088
rect 33376 36048 33382 36060
rect 33778 36048 33784 36060
rect 33836 36048 33842 36100
rect 33873 36091 33931 36097
rect 33873 36057 33885 36091
rect 33919 36088 33931 36091
rect 34882 36088 34888 36100
rect 33919 36060 34888 36088
rect 33919 36057 33931 36060
rect 33873 36051 33931 36057
rect 28350 35980 28356 36032
rect 28408 36020 28414 36032
rect 28997 36023 29055 36029
rect 28997 36020 29009 36023
rect 28408 35992 29009 36020
rect 28408 35980 28414 35992
rect 28997 35989 29009 35992
rect 29043 36020 29055 36023
rect 30650 36020 30656 36032
rect 29043 35992 30656 36020
rect 29043 35989 29055 35992
rect 28997 35983 29055 35989
rect 30650 35980 30656 35992
rect 30708 35980 30714 36032
rect 32490 35980 32496 36032
rect 32548 36020 32554 36032
rect 33888 36020 33916 36051
rect 34882 36048 34888 36060
rect 34940 36048 34946 36100
rect 35084 36088 35112 36119
rect 35986 36116 35992 36128
rect 36044 36116 36050 36168
rect 36556 36165 36584 36196
rect 36722 36184 36728 36196
rect 36780 36184 36786 36236
rect 37458 36184 37464 36236
rect 37516 36224 37522 36236
rect 37516 36196 37964 36224
rect 37516 36184 37522 36196
rect 36517 36159 36584 36165
rect 36517 36125 36529 36159
rect 36563 36128 36584 36159
rect 36633 36159 36691 36165
rect 36563 36125 36575 36128
rect 36517 36119 36575 36125
rect 36633 36125 36645 36159
rect 36679 36156 36691 36159
rect 37182 36156 37188 36168
rect 36679 36128 37188 36156
rect 36679 36125 36691 36128
rect 36633 36119 36691 36125
rect 37182 36116 37188 36128
rect 37240 36116 37246 36168
rect 37642 36156 37648 36168
rect 37603 36128 37648 36156
rect 37642 36116 37648 36128
rect 37700 36116 37706 36168
rect 37936 36165 37964 36196
rect 38125 36165 38153 36264
rect 40586 36252 40592 36304
rect 40644 36292 40650 36304
rect 42518 36292 42524 36304
rect 40644 36264 42524 36292
rect 40644 36252 40650 36264
rect 42518 36252 42524 36264
rect 42576 36292 42582 36304
rect 44361 36295 44419 36301
rect 44361 36292 44373 36295
rect 42576 36264 44373 36292
rect 42576 36252 42582 36264
rect 44361 36261 44373 36264
rect 44407 36261 44419 36295
rect 44361 36255 44419 36261
rect 44910 36252 44916 36304
rect 44968 36292 44974 36304
rect 46934 36292 46940 36304
rect 44968 36264 46940 36292
rect 44968 36252 44974 36264
rect 46934 36252 46940 36264
rect 46992 36292 46998 36304
rect 47581 36295 47639 36301
rect 47581 36292 47593 36295
rect 46992 36264 47593 36292
rect 46992 36252 46998 36264
rect 47581 36261 47593 36264
rect 47627 36261 47639 36295
rect 47581 36255 47639 36261
rect 47946 36252 47952 36304
rect 48004 36292 48010 36304
rect 50706 36292 50712 36304
rect 48004 36264 48268 36292
rect 48004 36252 48010 36264
rect 39942 36184 39948 36236
rect 40000 36224 40006 36236
rect 41141 36227 41199 36233
rect 40000 36196 41000 36224
rect 40000 36184 40006 36196
rect 37738 36159 37796 36165
rect 37738 36125 37750 36159
rect 37784 36125 37796 36159
rect 37738 36119 37796 36125
rect 37921 36159 37979 36165
rect 37921 36125 37933 36159
rect 37967 36125 37979 36159
rect 37921 36119 37979 36125
rect 38110 36159 38168 36165
rect 38110 36125 38122 36159
rect 38156 36125 38168 36159
rect 38110 36119 38168 36125
rect 37093 36091 37151 36097
rect 37093 36088 37105 36091
rect 35084 36060 37105 36088
rect 37093 36057 37105 36060
rect 37139 36057 37151 36091
rect 37093 36051 37151 36057
rect 32548 35992 33916 36020
rect 32548 35980 32554 35992
rect 34054 35980 34060 36032
rect 34112 36020 34118 36032
rect 34149 36023 34207 36029
rect 34149 36020 34161 36023
rect 34112 35992 34161 36020
rect 34112 35980 34118 35992
rect 34149 35989 34161 35992
rect 34195 35989 34207 36023
rect 34149 35983 34207 35989
rect 34606 35980 34612 36032
rect 34664 36020 34670 36032
rect 35253 36023 35311 36029
rect 35253 36020 35265 36023
rect 34664 35992 35265 36020
rect 34664 35980 34670 35992
rect 35253 35989 35265 35992
rect 35299 35989 35311 36023
rect 35253 35983 35311 35989
rect 35894 35980 35900 36032
rect 35952 36020 35958 36032
rect 36173 36023 36231 36029
rect 36173 36020 36185 36023
rect 35952 35992 36185 36020
rect 35952 35980 35958 35992
rect 36173 35989 36185 35992
rect 36219 35989 36231 36023
rect 36173 35983 36231 35989
rect 36265 36023 36323 36029
rect 36265 35989 36277 36023
rect 36311 36020 36323 36023
rect 36354 36020 36360 36032
rect 36311 35992 36360 36020
rect 36311 35989 36323 35992
rect 36265 35983 36323 35989
rect 36354 35980 36360 35992
rect 36412 35980 36418 36032
rect 37108 36020 37136 36051
rect 37550 36048 37556 36100
rect 37608 36088 37614 36100
rect 37752 36088 37780 36119
rect 38286 36116 38292 36168
rect 38344 36156 38350 36168
rect 38749 36159 38807 36165
rect 38749 36156 38761 36159
rect 38344 36128 38761 36156
rect 38344 36116 38350 36128
rect 38749 36125 38761 36128
rect 38795 36125 38807 36159
rect 38749 36119 38807 36125
rect 40037 36159 40095 36165
rect 40037 36125 40049 36159
rect 40083 36156 40095 36159
rect 40126 36156 40132 36168
rect 40083 36128 40132 36156
rect 40083 36125 40095 36128
rect 40037 36119 40095 36125
rect 40126 36116 40132 36128
rect 40184 36116 40190 36168
rect 40972 36165 41000 36196
rect 41141 36193 41153 36227
rect 41187 36224 41199 36227
rect 41506 36224 41512 36236
rect 41187 36196 41512 36224
rect 41187 36193 41199 36196
rect 41141 36187 41199 36193
rect 41506 36184 41512 36196
rect 41564 36184 41570 36236
rect 41782 36184 41788 36236
rect 41840 36224 41846 36236
rect 41969 36227 42027 36233
rect 41969 36224 41981 36227
rect 41840 36196 41981 36224
rect 41840 36184 41846 36196
rect 41969 36193 41981 36196
rect 42015 36193 42027 36227
rect 42886 36224 42892 36236
rect 42847 36196 42892 36224
rect 41969 36187 42027 36193
rect 42886 36184 42892 36196
rect 42944 36184 42950 36236
rect 42978 36184 42984 36236
rect 43036 36224 43042 36236
rect 44177 36227 44235 36233
rect 44177 36224 44189 36227
rect 43036 36196 44189 36224
rect 43036 36184 43042 36196
rect 44177 36193 44189 36196
rect 44223 36193 44235 36227
rect 44177 36187 44235 36193
rect 44269 36227 44327 36233
rect 44269 36193 44281 36227
rect 44315 36224 44327 36227
rect 45002 36224 45008 36236
rect 44315 36196 45008 36224
rect 44315 36193 44327 36196
rect 44269 36187 44327 36193
rect 45002 36184 45008 36196
rect 45060 36184 45066 36236
rect 45738 36224 45744 36236
rect 45699 36196 45744 36224
rect 45738 36184 45744 36196
rect 45796 36184 45802 36236
rect 46492 36196 48084 36224
rect 46492 36168 46520 36196
rect 40957 36159 41015 36165
rect 40957 36125 40969 36159
rect 41003 36156 41015 36159
rect 41874 36156 41880 36168
rect 41003 36128 41880 36156
rect 41003 36125 41015 36128
rect 40957 36119 41015 36125
rect 41874 36116 41880 36128
rect 41932 36116 41938 36168
rect 42245 36159 42303 36165
rect 42245 36125 42257 36159
rect 42291 36156 42303 36159
rect 42334 36156 42340 36168
rect 42291 36128 42340 36156
rect 42291 36125 42303 36128
rect 42245 36119 42303 36125
rect 42334 36116 42340 36128
rect 42392 36116 42398 36168
rect 42429 36159 42487 36165
rect 42429 36125 42441 36159
rect 42475 36125 42487 36159
rect 42429 36119 42487 36125
rect 38010 36088 38016 36100
rect 37608 36060 37780 36088
rect 37971 36060 38016 36088
rect 37608 36048 37614 36060
rect 38010 36048 38016 36060
rect 38068 36048 38074 36100
rect 41325 36091 41383 36097
rect 38212 36060 38516 36088
rect 38212 36020 38240 36060
rect 37108 35992 38240 36020
rect 38289 36023 38347 36029
rect 38289 35989 38301 36023
rect 38335 36020 38347 36023
rect 38378 36020 38384 36032
rect 38335 35992 38384 36020
rect 38335 35989 38347 35992
rect 38289 35983 38347 35989
rect 38378 35980 38384 35992
rect 38436 35980 38442 36032
rect 38488 36020 38516 36060
rect 41325 36057 41337 36091
rect 41371 36088 41383 36091
rect 42444 36088 42472 36119
rect 42610 36116 42616 36168
rect 42668 36156 42674 36168
rect 43073 36159 43131 36165
rect 43073 36156 43085 36159
rect 42668 36128 43085 36156
rect 42668 36116 42674 36128
rect 43073 36125 43085 36128
rect 43119 36125 43131 36159
rect 43073 36119 43131 36125
rect 43162 36116 43168 36168
rect 43220 36156 43226 36168
rect 43533 36159 43591 36165
rect 43220 36128 43265 36156
rect 43220 36116 43226 36128
rect 43533 36125 43545 36159
rect 43579 36156 43591 36159
rect 43993 36159 44051 36165
rect 43579 36128 43668 36156
rect 43579 36125 43591 36128
rect 43533 36119 43591 36125
rect 41371 36060 41736 36088
rect 41371 36057 41383 36060
rect 41325 36051 41383 36057
rect 38654 36020 38660 36032
rect 38488 35992 38660 36020
rect 38654 35980 38660 35992
rect 38712 36020 38718 36032
rect 39393 36023 39451 36029
rect 39393 36020 39405 36023
rect 38712 35992 39405 36020
rect 38712 35980 38718 35992
rect 39393 35989 39405 35992
rect 39439 36020 39451 36023
rect 40126 36020 40132 36032
rect 39439 35992 40132 36020
rect 39439 35989 39451 35992
rect 39393 35983 39451 35989
rect 40126 35980 40132 35992
rect 40184 35980 40190 36032
rect 40221 36023 40279 36029
rect 40221 35989 40233 36023
rect 40267 36020 40279 36023
rect 40678 36020 40684 36032
rect 40267 35992 40684 36020
rect 40267 35989 40279 35992
rect 40221 35983 40279 35989
rect 40678 35980 40684 35992
rect 40736 35980 40742 36032
rect 41708 36020 41736 36060
rect 42444 36060 42748 36088
rect 42444 36020 42472 36060
rect 42720 36032 42748 36060
rect 41708 35992 42472 36020
rect 42702 35980 42708 36032
rect 42760 36020 42766 36032
rect 43640 36020 43668 36128
rect 43993 36125 44005 36159
rect 44039 36156 44051 36159
rect 44039 36150 44220 36156
rect 44039 36128 44312 36150
rect 44039 36125 44051 36128
rect 43993 36119 44051 36125
rect 44192 36122 44312 36128
rect 44284 36088 44312 36122
rect 44450 36116 44456 36168
rect 44508 36156 44514 36168
rect 45557 36159 45615 36165
rect 45557 36156 45569 36159
rect 44508 36128 45569 36156
rect 44508 36116 44514 36128
rect 45557 36125 45569 36128
rect 45603 36125 45615 36159
rect 46474 36156 46480 36168
rect 46435 36128 46480 36156
rect 45557 36119 45615 36125
rect 46474 36116 46480 36128
rect 46532 36116 46538 36168
rect 46753 36159 46811 36165
rect 46753 36125 46765 36159
rect 46799 36156 46811 36159
rect 46842 36156 46848 36168
rect 46799 36128 46848 36156
rect 46799 36125 46811 36128
rect 46753 36119 46811 36125
rect 44910 36088 44916 36100
rect 44284 36060 44916 36088
rect 44910 36048 44916 36060
rect 44968 36048 44974 36100
rect 45649 36091 45707 36097
rect 45649 36057 45661 36091
rect 45695 36088 45707 36091
rect 46768 36088 46796 36119
rect 46842 36116 46848 36128
rect 46900 36116 46906 36168
rect 47394 36156 47400 36168
rect 47355 36128 47400 36156
rect 47394 36116 47400 36128
rect 47452 36116 47458 36168
rect 47578 36156 47584 36168
rect 47539 36128 47584 36156
rect 47578 36116 47584 36128
rect 47636 36116 47642 36168
rect 48056 36165 48084 36196
rect 48240 36165 48268 36264
rect 50448 36264 50712 36292
rect 48682 36184 48688 36236
rect 48740 36224 48746 36236
rect 48869 36227 48927 36233
rect 48869 36224 48881 36227
rect 48740 36196 48881 36224
rect 48740 36184 48746 36196
rect 48869 36193 48881 36196
rect 48915 36224 48927 36227
rect 49694 36224 49700 36236
rect 48915 36196 49700 36224
rect 48915 36193 48927 36196
rect 48869 36187 48927 36193
rect 49694 36184 49700 36196
rect 49752 36224 49758 36236
rect 50448 36224 50476 36264
rect 50706 36252 50712 36264
rect 50764 36252 50770 36304
rect 53101 36295 53159 36301
rect 53101 36261 53113 36295
rect 53147 36261 53159 36295
rect 53101 36255 53159 36261
rect 50982 36224 50988 36236
rect 49752 36196 50476 36224
rect 49752 36184 49758 36196
rect 48041 36159 48099 36165
rect 48041 36125 48053 36159
rect 48087 36125 48099 36159
rect 48041 36119 48099 36125
rect 48225 36159 48283 36165
rect 48225 36125 48237 36159
rect 48271 36125 48283 36159
rect 49050 36156 49056 36168
rect 49011 36128 49056 36156
rect 48225 36119 48283 36125
rect 49050 36116 49056 36128
rect 49108 36116 49114 36168
rect 50338 36156 50344 36168
rect 50299 36128 50344 36156
rect 50338 36116 50344 36128
rect 50396 36116 50402 36168
rect 50448 36165 50476 36196
rect 50632 36196 50988 36224
rect 50632 36168 50660 36196
rect 50982 36184 50988 36196
rect 51040 36184 51046 36236
rect 52822 36224 52828 36236
rect 52783 36196 52828 36224
rect 52822 36184 52828 36196
rect 52880 36184 52886 36236
rect 53116 36224 53144 36255
rect 53929 36227 53987 36233
rect 53929 36224 53941 36227
rect 53116 36196 53941 36224
rect 53929 36193 53941 36196
rect 53975 36193 53987 36227
rect 53929 36187 53987 36193
rect 50434 36159 50492 36165
rect 50434 36125 50446 36159
rect 50480 36125 50492 36159
rect 50434 36119 50492 36125
rect 50614 36116 50620 36168
rect 50672 36156 50678 36168
rect 50890 36165 50896 36168
rect 50847 36159 50896 36165
rect 50672 36128 50765 36156
rect 50672 36116 50678 36128
rect 50847 36125 50859 36159
rect 50893 36125 50896 36159
rect 50847 36119 50896 36125
rect 50890 36116 50896 36119
rect 50948 36156 50954 36168
rect 51258 36156 51264 36168
rect 50948 36128 51264 36156
rect 50948 36116 50954 36128
rect 51258 36116 51264 36128
rect 51316 36116 51322 36168
rect 52730 36156 52736 36168
rect 52691 36128 52736 36156
rect 52730 36116 52736 36128
rect 52788 36116 52794 36168
rect 53282 36116 53288 36168
rect 53340 36156 53346 36168
rect 53650 36156 53656 36168
rect 53340 36128 53656 36156
rect 53340 36116 53346 36128
rect 53650 36116 53656 36128
rect 53708 36156 53714 36168
rect 54021 36159 54079 36165
rect 54021 36156 54033 36159
rect 53708 36128 54033 36156
rect 53708 36116 53714 36128
rect 54021 36125 54033 36128
rect 54067 36125 54079 36159
rect 54021 36119 54079 36125
rect 55122 36116 55128 36168
rect 55180 36156 55186 36168
rect 55861 36159 55919 36165
rect 55861 36156 55873 36159
rect 55180 36128 55873 36156
rect 55180 36116 55186 36128
rect 55861 36125 55873 36128
rect 55907 36125 55919 36159
rect 56134 36156 56140 36168
rect 56095 36128 56140 36156
rect 55861 36119 55919 36125
rect 56134 36116 56140 36128
rect 56192 36116 56198 36168
rect 57422 36156 57428 36168
rect 57383 36128 57428 36156
rect 57422 36116 57428 36128
rect 57480 36116 57486 36168
rect 57698 36156 57704 36168
rect 57659 36128 57704 36156
rect 57698 36116 57704 36128
rect 57756 36116 57762 36168
rect 45695 36060 46796 36088
rect 46937 36091 46995 36097
rect 45695 36057 45707 36060
rect 45649 36051 45707 36057
rect 46937 36057 46949 36091
rect 46983 36088 46995 36091
rect 48406 36088 48412 36100
rect 46983 36060 48412 36088
rect 46983 36057 46995 36060
rect 46937 36051 46995 36057
rect 48406 36048 48412 36060
rect 48464 36048 48470 36100
rect 50062 36048 50068 36100
rect 50120 36088 50126 36100
rect 50709 36091 50767 36097
rect 50709 36088 50721 36091
rect 50120 36060 50721 36088
rect 50120 36048 50126 36060
rect 50709 36057 50721 36060
rect 50755 36057 50767 36091
rect 50709 36051 50767 36057
rect 44266 36020 44272 36032
rect 42760 35992 44272 36020
rect 42760 35980 42766 35992
rect 44266 35980 44272 35992
rect 44324 35980 44330 36032
rect 45186 36020 45192 36032
rect 45147 35992 45192 36020
rect 45186 35980 45192 35992
rect 45244 35980 45250 36032
rect 46566 36020 46572 36032
rect 46527 35992 46572 36020
rect 46566 35980 46572 35992
rect 46624 36020 46630 36032
rect 47946 36020 47952 36032
rect 46624 35992 47952 36020
rect 46624 35980 46630 35992
rect 47946 35980 47952 35992
rect 48004 35980 48010 36032
rect 48130 36020 48136 36032
rect 48091 35992 48136 36020
rect 48130 35980 48136 35992
rect 48188 35980 48194 36032
rect 48498 35980 48504 36032
rect 48556 36020 48562 36032
rect 49237 36023 49295 36029
rect 49237 36020 49249 36023
rect 48556 35992 49249 36020
rect 48556 35980 48562 35992
rect 49237 35989 49249 35992
rect 49283 36020 49295 36023
rect 49326 36020 49332 36032
rect 49283 35992 49332 36020
rect 49283 35989 49295 35992
rect 49237 35983 49295 35989
rect 49326 35980 49332 35992
rect 49384 35980 49390 36032
rect 50798 35980 50804 36032
rect 50856 36020 50862 36032
rect 50985 36023 51043 36029
rect 50985 36020 50997 36023
rect 50856 35992 50997 36020
rect 50856 35980 50862 35992
rect 50985 35989 50997 35992
rect 51031 35989 51043 36023
rect 51626 36020 51632 36032
rect 51587 35992 51632 36020
rect 50985 35983 51043 35989
rect 51626 35980 51632 35992
rect 51684 35980 51690 36032
rect 52086 35980 52092 36032
rect 52144 36020 52150 36032
rect 54294 36020 54300 36032
rect 52144 35992 54300 36020
rect 52144 35980 52150 35992
rect 54294 35980 54300 35992
rect 54352 36020 54358 36032
rect 54662 36020 54668 36032
rect 54352 35992 54668 36020
rect 54352 35980 54358 35992
rect 54662 35980 54668 35992
rect 54720 35980 54726 36032
rect 54846 36020 54852 36032
rect 54807 35992 54852 36020
rect 54846 35980 54852 35992
rect 54904 35980 54910 36032
rect 55214 35980 55220 36032
rect 55272 36020 55278 36032
rect 55493 36023 55551 36029
rect 55493 36020 55505 36023
rect 55272 35992 55505 36020
rect 55272 35980 55278 35992
rect 55493 35989 55505 35992
rect 55539 35989 55551 36023
rect 55493 35983 55551 35989
rect 56870 35980 56876 36032
rect 56928 36020 56934 36032
rect 57057 36023 57115 36029
rect 57057 36020 57069 36023
rect 56928 35992 57069 36020
rect 56928 35980 56934 35992
rect 57057 35989 57069 35992
rect 57103 35989 57115 36023
rect 57057 35983 57115 35989
rect 1104 35930 58880 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 58880 35930
rect 1104 35856 58880 35878
rect 29089 35819 29147 35825
rect 29089 35785 29101 35819
rect 29135 35816 29147 35819
rect 29454 35816 29460 35828
rect 29135 35788 29460 35816
rect 29135 35785 29147 35788
rect 29089 35779 29147 35785
rect 29454 35776 29460 35788
rect 29512 35816 29518 35828
rect 30282 35816 30288 35828
rect 29512 35788 30288 35816
rect 29512 35776 29518 35788
rect 30282 35776 30288 35788
rect 30340 35816 30346 35828
rect 31662 35816 31668 35828
rect 30340 35788 31668 35816
rect 30340 35776 30346 35788
rect 31662 35776 31668 35788
rect 31720 35776 31726 35828
rect 32677 35819 32735 35825
rect 32677 35785 32689 35819
rect 32723 35816 32735 35819
rect 32723 35788 34376 35816
rect 32723 35785 32735 35788
rect 32677 35779 32735 35785
rect 28902 35708 28908 35760
rect 28960 35748 28966 35760
rect 30377 35751 30435 35757
rect 28960 35720 30236 35748
rect 28960 35708 28966 35720
rect 29012 35689 29040 35720
rect 28997 35683 29055 35689
rect 28997 35649 29009 35683
rect 29043 35649 29055 35683
rect 28997 35643 29055 35649
rect 29178 35640 29184 35692
rect 29236 35680 29242 35692
rect 29273 35683 29331 35689
rect 29273 35680 29285 35683
rect 29236 35652 29285 35680
rect 29236 35640 29242 35652
rect 29273 35649 29285 35652
rect 29319 35649 29331 35683
rect 30098 35680 30104 35692
rect 30059 35652 30104 35680
rect 29273 35643 29331 35649
rect 29288 35612 29316 35643
rect 30098 35640 30104 35652
rect 30156 35640 30162 35692
rect 30208 35680 30236 35720
rect 30377 35717 30389 35751
rect 30423 35748 30435 35751
rect 30558 35748 30564 35760
rect 30423 35720 30564 35748
rect 30423 35717 30435 35720
rect 30377 35711 30435 35717
rect 30558 35708 30564 35720
rect 30616 35748 30622 35760
rect 31294 35748 31300 35760
rect 30616 35720 31300 35748
rect 30616 35708 30622 35720
rect 31294 35708 31300 35720
rect 31352 35708 31358 35760
rect 31202 35680 31208 35692
rect 30208 35652 31208 35680
rect 31202 35640 31208 35652
rect 31260 35640 31266 35692
rect 31386 35680 31392 35692
rect 31347 35652 31392 35680
rect 31386 35640 31392 35652
rect 31444 35640 31450 35692
rect 31757 35683 31815 35689
rect 31757 35649 31769 35683
rect 31803 35680 31815 35683
rect 32692 35680 32720 35779
rect 33594 35748 33600 35760
rect 33555 35720 33600 35748
rect 33594 35708 33600 35720
rect 33652 35708 33658 35760
rect 33318 35680 33324 35692
rect 31803 35652 32720 35680
rect 32784 35652 33324 35680
rect 31803 35649 31815 35652
rect 31757 35643 31815 35649
rect 32493 35615 32551 35621
rect 29288 35584 31754 35612
rect 29270 35544 29276 35556
rect 29231 35516 29276 35544
rect 29270 35504 29276 35516
rect 29328 35504 29334 35556
rect 31726 35544 31754 35584
rect 32493 35581 32505 35615
rect 32539 35612 32551 35615
rect 32784 35612 32812 35652
rect 33318 35640 33324 35652
rect 33376 35640 33382 35692
rect 34054 35640 34060 35692
rect 34112 35640 34118 35692
rect 34348 35680 34376 35788
rect 34698 35776 34704 35828
rect 34756 35816 34762 35828
rect 35437 35819 35495 35825
rect 35437 35816 35449 35819
rect 34756 35788 35449 35816
rect 34756 35776 34762 35788
rect 35437 35785 35449 35788
rect 35483 35816 35495 35819
rect 35710 35816 35716 35828
rect 35483 35788 35716 35816
rect 35483 35785 35495 35788
rect 35437 35779 35495 35785
rect 35710 35776 35716 35788
rect 35768 35776 35774 35828
rect 35805 35819 35863 35825
rect 35805 35785 35817 35819
rect 35851 35785 35863 35819
rect 35805 35779 35863 35785
rect 34882 35708 34888 35760
rect 34940 35748 34946 35760
rect 35820 35748 35848 35779
rect 37458 35776 37464 35828
rect 37516 35816 37522 35828
rect 38930 35816 38936 35828
rect 37516 35788 38936 35816
rect 37516 35776 37522 35788
rect 38930 35776 38936 35788
rect 38988 35776 38994 35828
rect 41414 35776 41420 35828
rect 41472 35816 41478 35828
rect 41509 35819 41567 35825
rect 41509 35816 41521 35819
rect 41472 35788 41521 35816
rect 41472 35776 41478 35788
rect 41509 35785 41521 35788
rect 41555 35785 41567 35819
rect 42702 35816 42708 35828
rect 42663 35788 42708 35816
rect 41509 35779 41567 35785
rect 38289 35751 38347 35757
rect 38289 35748 38301 35751
rect 34940 35720 35664 35748
rect 35820 35720 38301 35748
rect 34940 35708 34946 35720
rect 35636 35680 35664 35720
rect 38289 35717 38301 35720
rect 38335 35717 38347 35751
rect 38289 35711 38347 35717
rect 38473 35751 38531 35757
rect 38473 35717 38485 35751
rect 38519 35748 38531 35751
rect 38838 35748 38844 35760
rect 38519 35720 38844 35748
rect 38519 35717 38531 35720
rect 38473 35711 38531 35717
rect 38838 35708 38844 35720
rect 38896 35708 38902 35760
rect 41524 35748 41552 35779
rect 42702 35776 42708 35788
rect 42760 35776 42766 35828
rect 43070 35816 43076 35828
rect 43031 35788 43076 35816
rect 43070 35776 43076 35788
rect 43128 35776 43134 35828
rect 44177 35819 44235 35825
rect 44177 35785 44189 35819
rect 44223 35816 44235 35819
rect 44450 35816 44456 35828
rect 44223 35788 44456 35816
rect 44223 35785 44235 35788
rect 44177 35779 44235 35785
rect 44450 35776 44456 35788
rect 44508 35776 44514 35828
rect 45005 35819 45063 35825
rect 45005 35785 45017 35819
rect 45051 35816 45063 35819
rect 45373 35819 45431 35825
rect 45051 35788 45324 35816
rect 45051 35785 45063 35788
rect 45005 35779 45063 35785
rect 41524 35720 42288 35748
rect 36265 35683 36323 35689
rect 36265 35680 36277 35683
rect 34348 35652 35572 35680
rect 35636 35652 36277 35680
rect 32539 35584 32812 35612
rect 32539 35581 32551 35584
rect 32493 35575 32551 35581
rect 32858 35572 32864 35624
rect 32916 35612 32922 35624
rect 34149 35615 34207 35621
rect 34149 35612 34161 35615
rect 32916 35584 32961 35612
rect 33060 35584 34161 35612
rect 32916 35572 32922 35584
rect 32766 35544 32772 35556
rect 31726 35516 32772 35544
rect 32766 35504 32772 35516
rect 32824 35504 32830 35556
rect 32306 35476 32312 35488
rect 32267 35448 32312 35476
rect 32306 35436 32312 35448
rect 32364 35436 32370 35488
rect 32398 35436 32404 35488
rect 32456 35476 32462 35488
rect 32876 35476 32904 35572
rect 32950 35504 32956 35556
rect 33008 35544 33014 35556
rect 33060 35544 33088 35584
rect 34149 35581 34161 35584
rect 34195 35581 34207 35615
rect 34149 35575 34207 35581
rect 35253 35615 35311 35621
rect 35253 35581 35265 35615
rect 35299 35581 35311 35615
rect 35253 35575 35311 35581
rect 33008 35516 33088 35544
rect 35268 35544 35296 35575
rect 35342 35572 35348 35624
rect 35400 35612 35406 35624
rect 35400 35584 35445 35612
rect 35400 35572 35406 35584
rect 35434 35544 35440 35556
rect 35268 35516 35440 35544
rect 33008 35504 33014 35516
rect 35434 35504 35440 35516
rect 35492 35504 35498 35556
rect 35544 35544 35572 35652
rect 36265 35649 36277 35652
rect 36311 35680 36323 35683
rect 36538 35680 36544 35692
rect 36311 35652 36544 35680
rect 36311 35649 36323 35652
rect 36265 35643 36323 35649
rect 36538 35640 36544 35652
rect 36596 35640 36602 35692
rect 37458 35680 37464 35692
rect 37419 35652 37464 35680
rect 37458 35640 37464 35652
rect 37516 35640 37522 35692
rect 37550 35640 37556 35692
rect 37608 35680 37614 35692
rect 37608 35652 37653 35680
rect 37608 35640 37614 35652
rect 37734 35640 37740 35692
rect 37792 35680 37798 35692
rect 38562 35680 38568 35692
rect 37792 35652 37837 35680
rect 38523 35652 38568 35680
rect 37792 35640 37798 35652
rect 38562 35640 38568 35652
rect 38620 35640 38626 35692
rect 39206 35680 39212 35692
rect 39167 35652 39212 35680
rect 39206 35640 39212 35652
rect 39264 35640 39270 35692
rect 40221 35683 40279 35689
rect 40221 35649 40233 35683
rect 40267 35680 40279 35683
rect 40862 35680 40868 35692
rect 40267 35652 40868 35680
rect 40267 35649 40279 35652
rect 40221 35643 40279 35649
rect 40862 35640 40868 35652
rect 40920 35640 40926 35692
rect 41414 35640 41420 35692
rect 41472 35680 41478 35692
rect 41601 35683 41659 35689
rect 41472 35652 41517 35680
rect 41472 35640 41478 35652
rect 41601 35649 41613 35683
rect 41647 35680 41659 35683
rect 41874 35680 41880 35692
rect 41647 35652 41880 35680
rect 41647 35649 41659 35652
rect 41601 35643 41659 35649
rect 41874 35640 41880 35652
rect 41932 35640 41938 35692
rect 42260 35680 42288 35720
rect 42610 35680 42616 35692
rect 42260 35652 42616 35680
rect 42610 35640 42616 35652
rect 42668 35640 42674 35692
rect 42889 35683 42947 35689
rect 42889 35649 42901 35683
rect 42935 35680 42947 35683
rect 43162 35680 43168 35692
rect 42935 35652 43168 35680
rect 42935 35649 42947 35652
rect 42889 35643 42947 35649
rect 43162 35640 43168 35652
rect 43220 35640 43226 35692
rect 44082 35680 44088 35692
rect 44043 35652 44088 35680
rect 44082 35640 44088 35652
rect 44140 35640 44146 35692
rect 44174 35640 44180 35692
rect 44232 35680 44238 35692
rect 44913 35683 44971 35689
rect 44913 35680 44925 35683
rect 44232 35652 44925 35680
rect 44232 35640 44238 35652
rect 44913 35649 44925 35652
rect 44959 35649 44971 35683
rect 45186 35680 45192 35692
rect 45147 35652 45192 35680
rect 44913 35643 44971 35649
rect 45186 35640 45192 35652
rect 45244 35640 45250 35692
rect 45296 35680 45324 35788
rect 45373 35785 45385 35819
rect 45419 35816 45431 35819
rect 45738 35816 45744 35828
rect 45419 35788 45744 35816
rect 45419 35785 45431 35788
rect 45373 35779 45431 35785
rect 45738 35776 45744 35788
rect 45796 35776 45802 35828
rect 48700 35788 50752 35816
rect 46106 35708 46112 35760
rect 46164 35748 46170 35760
rect 46164 35720 46428 35748
rect 46164 35708 46170 35720
rect 45922 35680 45928 35692
rect 45296 35652 45928 35680
rect 45922 35640 45928 35652
rect 45980 35680 45986 35692
rect 46017 35683 46075 35689
rect 46017 35680 46029 35683
rect 45980 35652 46029 35680
rect 45980 35640 45986 35652
rect 46017 35649 46029 35652
rect 46063 35649 46075 35683
rect 46198 35680 46204 35692
rect 46159 35652 46204 35680
rect 46017 35643 46075 35649
rect 46198 35640 46204 35652
rect 46256 35640 46262 35692
rect 46400 35689 46428 35720
rect 46293 35683 46351 35689
rect 46293 35649 46305 35683
rect 46339 35649 46351 35683
rect 46293 35643 46351 35649
rect 46385 35683 46443 35689
rect 46385 35649 46397 35683
rect 46431 35649 46443 35683
rect 46385 35643 46443 35649
rect 47213 35683 47271 35689
rect 47213 35649 47225 35683
rect 47259 35680 47271 35683
rect 47946 35680 47952 35692
rect 47259 35652 47952 35680
rect 47259 35649 47271 35652
rect 47213 35643 47271 35649
rect 39117 35615 39175 35621
rect 39117 35612 39129 35615
rect 38304 35584 39129 35612
rect 37182 35544 37188 35556
rect 35544 35516 37188 35544
rect 37182 35504 37188 35516
rect 37240 35504 37246 35556
rect 37642 35504 37648 35556
rect 37700 35544 37706 35556
rect 38304 35553 38332 35584
rect 39117 35581 39129 35584
rect 39163 35581 39175 35615
rect 40129 35615 40187 35621
rect 40129 35612 40141 35615
rect 39117 35575 39175 35581
rect 39592 35584 40141 35612
rect 39592 35553 39620 35584
rect 40129 35581 40141 35584
rect 40175 35581 40187 35615
rect 46308 35612 46336 35643
rect 47946 35640 47952 35652
rect 48004 35640 48010 35692
rect 47118 35612 47124 35624
rect 40129 35575 40187 35581
rect 41386 35584 47124 35612
rect 37737 35547 37795 35553
rect 37737 35544 37749 35547
rect 37700 35516 37749 35544
rect 37700 35504 37706 35516
rect 37737 35513 37749 35516
rect 37783 35513 37795 35547
rect 37737 35507 37795 35513
rect 38289 35547 38347 35553
rect 38289 35513 38301 35547
rect 38335 35513 38347 35547
rect 38289 35507 38347 35513
rect 39577 35547 39635 35553
rect 39577 35513 39589 35547
rect 39623 35513 39635 35547
rect 39577 35507 39635 35513
rect 40589 35547 40647 35553
rect 40589 35513 40601 35547
rect 40635 35544 40647 35547
rect 40954 35544 40960 35556
rect 40635 35516 40960 35544
rect 40635 35513 40647 35516
rect 40589 35507 40647 35513
rect 40954 35504 40960 35516
rect 41012 35504 41018 35556
rect 32456 35448 32904 35476
rect 32456 35436 32462 35448
rect 36170 35436 36176 35488
rect 36228 35476 36234 35488
rect 36357 35479 36415 35485
rect 36357 35476 36369 35479
rect 36228 35448 36369 35476
rect 36228 35436 36234 35448
rect 36357 35445 36369 35448
rect 36403 35476 36415 35479
rect 41386 35476 41414 35584
rect 47118 35572 47124 35584
rect 47176 35572 47182 35624
rect 47302 35572 47308 35624
rect 47360 35612 47366 35624
rect 48041 35615 48099 35621
rect 48041 35612 48053 35615
rect 47360 35584 48053 35612
rect 47360 35572 47366 35584
rect 48041 35581 48053 35584
rect 48087 35612 48099 35615
rect 48700 35612 48728 35788
rect 49881 35751 49939 35757
rect 49881 35717 49893 35751
rect 49927 35748 49939 35751
rect 50614 35748 50620 35760
rect 49927 35720 50476 35748
rect 50575 35720 50620 35748
rect 49927 35717 49939 35720
rect 49881 35711 49939 35717
rect 48774 35640 48780 35692
rect 48832 35680 48838 35692
rect 49145 35683 49203 35689
rect 49145 35680 49157 35683
rect 48832 35652 48877 35680
rect 49068 35652 49157 35680
rect 48832 35640 48838 35652
rect 48087 35584 48728 35612
rect 48087 35581 48099 35584
rect 48041 35575 48099 35581
rect 48866 35572 48872 35624
rect 48924 35612 48930 35624
rect 48961 35615 49019 35621
rect 48961 35612 48973 35615
rect 48924 35584 48973 35612
rect 48924 35572 48930 35584
rect 48961 35581 48973 35584
rect 49007 35581 49019 35615
rect 48961 35575 49019 35581
rect 44082 35504 44088 35556
rect 44140 35544 44146 35556
rect 46198 35544 46204 35556
rect 44140 35516 46204 35544
rect 44140 35504 44146 35516
rect 46198 35504 46204 35516
rect 46256 35504 46262 35556
rect 48314 35544 48320 35556
rect 48275 35516 48320 35544
rect 48314 35504 48320 35516
rect 48372 35504 48378 35556
rect 48682 35504 48688 35556
rect 48740 35544 48746 35556
rect 49068 35544 49096 35652
rect 49145 35649 49157 35652
rect 49191 35649 49203 35683
rect 49145 35643 49203 35649
rect 50246 35640 50252 35692
rect 50304 35680 50310 35692
rect 50448 35689 50476 35720
rect 50614 35708 50620 35720
rect 50672 35708 50678 35760
rect 50724 35748 50752 35788
rect 50982 35776 50988 35828
rect 51040 35816 51046 35828
rect 52270 35816 52276 35828
rect 51040 35788 52276 35816
rect 51040 35776 51046 35788
rect 52270 35776 52276 35788
rect 52328 35816 52334 35828
rect 56321 35819 56379 35825
rect 52328 35788 54984 35816
rect 52328 35776 52334 35788
rect 50724 35720 51074 35748
rect 50341 35683 50399 35689
rect 50341 35680 50353 35683
rect 50304 35652 50353 35680
rect 50304 35640 50310 35652
rect 50341 35649 50353 35652
rect 50387 35649 50399 35683
rect 50341 35643 50399 35649
rect 50434 35683 50492 35689
rect 50434 35649 50446 35683
rect 50480 35680 50492 35683
rect 50706 35680 50712 35692
rect 50480 35652 50568 35680
rect 50667 35652 50712 35680
rect 50480 35649 50492 35652
rect 50434 35643 50492 35649
rect 48740 35516 49096 35544
rect 49145 35547 49203 35553
rect 48740 35504 48746 35516
rect 49145 35513 49157 35547
rect 49191 35544 49203 35547
rect 49970 35544 49976 35556
rect 49191 35516 49976 35544
rect 49191 35513 49203 35516
rect 49145 35507 49203 35513
rect 49970 35504 49976 35516
rect 50028 35504 50034 35556
rect 36403 35448 41414 35476
rect 43625 35479 43683 35485
rect 36403 35445 36415 35448
rect 36357 35439 36415 35445
rect 43625 35445 43637 35479
rect 43671 35476 43683 35479
rect 45462 35476 45468 35488
rect 43671 35448 45468 35476
rect 43671 35445 43683 35448
rect 43625 35439 43683 35445
rect 45462 35436 45468 35448
rect 45520 35436 45526 35488
rect 46658 35476 46664 35488
rect 46619 35448 46664 35476
rect 46658 35436 46664 35448
rect 46716 35436 46722 35488
rect 50540 35476 50568 35652
rect 50706 35640 50712 35652
rect 50764 35640 50770 35692
rect 50847 35683 50905 35689
rect 50847 35680 50859 35683
rect 50821 35649 50859 35680
rect 50893 35649 50905 35683
rect 51046 35680 51074 35720
rect 54662 35708 54668 35760
rect 54720 35748 54726 35760
rect 54757 35751 54815 35757
rect 54757 35748 54769 35751
rect 54720 35720 54769 35748
rect 54720 35708 54726 35720
rect 54757 35717 54769 35720
rect 54803 35717 54815 35751
rect 54757 35711 54815 35717
rect 51629 35683 51687 35689
rect 51629 35680 51641 35683
rect 51046 35652 51641 35680
rect 50821 35643 50905 35649
rect 51629 35649 51641 35652
rect 51675 35649 51687 35683
rect 51629 35643 51687 35649
rect 50614 35572 50620 35624
rect 50672 35612 50678 35624
rect 50821 35612 50849 35643
rect 52730 35640 52736 35692
rect 52788 35680 52794 35692
rect 53193 35683 53251 35689
rect 53193 35680 53205 35683
rect 52788 35652 53205 35680
rect 52788 35640 52794 35652
rect 53193 35649 53205 35652
rect 53239 35649 53251 35683
rect 53193 35643 53251 35649
rect 53650 35640 53656 35692
rect 53708 35680 53714 35692
rect 54481 35683 54539 35689
rect 54481 35680 54493 35683
rect 53708 35652 54493 35680
rect 53708 35640 53714 35652
rect 54481 35649 54493 35652
rect 54527 35649 54539 35683
rect 54481 35643 54539 35649
rect 54570 35640 54576 35692
rect 54628 35680 54634 35692
rect 54956 35689 54984 35788
rect 56321 35785 56333 35819
rect 56367 35816 56379 35819
rect 57422 35816 57428 35828
rect 56367 35788 57428 35816
rect 56367 35785 56379 35788
rect 56321 35779 56379 35785
rect 57422 35776 57428 35788
rect 57480 35776 57486 35828
rect 56686 35708 56692 35760
rect 56744 35748 56750 35760
rect 56781 35751 56839 35757
rect 56781 35748 56793 35751
rect 56744 35720 56793 35748
rect 56744 35708 56750 35720
rect 56781 35717 56793 35720
rect 56827 35717 56839 35751
rect 57330 35748 57336 35760
rect 57291 35720 57336 35748
rect 56781 35711 56839 35717
rect 57330 35708 57336 35720
rect 57388 35708 57394 35760
rect 54849 35683 54907 35689
rect 54849 35680 54861 35683
rect 54628 35652 54721 35680
rect 54772 35652 54861 35680
rect 54628 35640 54634 35652
rect 50672 35584 50849 35612
rect 50672 35572 50678 35584
rect 50821 35544 50849 35584
rect 51537 35615 51595 35621
rect 51537 35581 51549 35615
rect 51583 35581 51595 35615
rect 53101 35615 53159 35621
rect 53101 35612 53113 35615
rect 51537 35575 51595 35581
rect 52012 35584 53113 35612
rect 50890 35544 50896 35556
rect 50821 35516 50896 35544
rect 50890 35504 50896 35516
rect 50948 35504 50954 35556
rect 50985 35547 51043 35553
rect 50985 35513 50997 35547
rect 51031 35544 51043 35547
rect 51552 35544 51580 35575
rect 52012 35553 52040 35584
rect 53101 35581 53113 35584
rect 53147 35581 53159 35615
rect 53101 35575 53159 35581
rect 53466 35572 53472 35624
rect 53524 35612 53530 35624
rect 53929 35615 53987 35621
rect 53929 35612 53941 35615
rect 53524 35584 53941 35612
rect 53524 35572 53530 35584
rect 53929 35581 53941 35584
rect 53975 35581 53987 35615
rect 53929 35575 53987 35581
rect 51031 35516 51580 35544
rect 51997 35547 52055 35553
rect 51031 35513 51043 35516
rect 50985 35507 51043 35513
rect 51997 35513 52009 35547
rect 52043 35513 52055 35547
rect 51997 35507 52055 35513
rect 51902 35476 51908 35488
rect 50540 35448 51908 35476
rect 51902 35436 51908 35448
rect 51960 35436 51966 35488
rect 54680 35476 54708 35652
rect 54772 35624 54800 35652
rect 54849 35649 54861 35652
rect 54895 35649 54907 35683
rect 54849 35643 54907 35649
rect 54946 35683 55004 35689
rect 54946 35649 54958 35683
rect 54992 35649 55004 35683
rect 54946 35643 55004 35649
rect 55953 35683 56011 35689
rect 55953 35649 55965 35683
rect 55999 35680 56011 35683
rect 56134 35680 56140 35692
rect 55999 35652 56140 35680
rect 55999 35649 56011 35652
rect 55953 35643 56011 35649
rect 56134 35640 56140 35652
rect 56192 35640 56198 35692
rect 54754 35572 54760 35624
rect 54812 35572 54818 35624
rect 55861 35615 55919 35621
rect 55861 35581 55873 35615
rect 55907 35581 55919 35615
rect 55861 35575 55919 35581
rect 55125 35547 55183 35553
rect 55125 35513 55137 35547
rect 55171 35544 55183 35547
rect 55876 35544 55904 35575
rect 55171 35516 55904 35544
rect 55171 35513 55183 35516
rect 55125 35507 55183 35513
rect 55398 35476 55404 35488
rect 54680 35448 55404 35476
rect 55398 35436 55404 35448
rect 55456 35436 55462 35488
rect 57698 35436 57704 35488
rect 57756 35476 57762 35488
rect 58069 35479 58127 35485
rect 58069 35476 58081 35479
rect 57756 35448 58081 35476
rect 57756 35436 57762 35448
rect 58069 35445 58081 35448
rect 58115 35445 58127 35479
rect 58069 35439 58127 35445
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 29181 35275 29239 35281
rect 29181 35241 29193 35275
rect 29227 35272 29239 35275
rect 30098 35272 30104 35284
rect 29227 35244 30104 35272
rect 29227 35241 29239 35244
rect 29181 35235 29239 35241
rect 30098 35232 30104 35244
rect 30156 35232 30162 35284
rect 30653 35275 30711 35281
rect 30653 35241 30665 35275
rect 30699 35272 30711 35275
rect 31202 35272 31208 35284
rect 30699 35244 31208 35272
rect 30699 35241 30711 35244
rect 30653 35235 30711 35241
rect 31202 35232 31208 35244
rect 31260 35232 31266 35284
rect 32030 35232 32036 35284
rect 32088 35272 32094 35284
rect 33413 35275 33471 35281
rect 32088 35244 32904 35272
rect 32088 35232 32094 35244
rect 32766 35204 32772 35216
rect 32727 35176 32772 35204
rect 32766 35164 32772 35176
rect 32824 35164 32830 35216
rect 32876 35204 32904 35244
rect 33413 35241 33425 35275
rect 33459 35272 33471 35275
rect 33502 35272 33508 35284
rect 33459 35244 33508 35272
rect 33459 35241 33471 35244
rect 33413 35235 33471 35241
rect 33502 35232 33508 35244
rect 33560 35232 33566 35284
rect 33870 35232 33876 35284
rect 33928 35272 33934 35284
rect 34885 35275 34943 35281
rect 34885 35272 34897 35275
rect 33928 35244 34897 35272
rect 33928 35232 33934 35244
rect 34885 35241 34897 35244
rect 34931 35241 34943 35275
rect 35434 35272 35440 35284
rect 35395 35244 35440 35272
rect 34885 35235 34943 35241
rect 35434 35232 35440 35244
rect 35492 35232 35498 35284
rect 37734 35272 37740 35284
rect 35820 35244 37740 35272
rect 33888 35204 33916 35232
rect 32876 35176 33916 35204
rect 33962 35164 33968 35216
rect 34020 35204 34026 35216
rect 34241 35207 34299 35213
rect 34241 35204 34253 35207
rect 34020 35176 34253 35204
rect 34020 35164 34026 35176
rect 34241 35173 34253 35176
rect 34287 35204 34299 35207
rect 35820 35204 35848 35244
rect 37734 35232 37740 35244
rect 37792 35232 37798 35284
rect 37826 35232 37832 35284
rect 37884 35272 37890 35284
rect 39301 35275 39359 35281
rect 39301 35272 39313 35275
rect 37884 35244 39313 35272
rect 37884 35232 37890 35244
rect 39301 35241 39313 35244
rect 39347 35241 39359 35275
rect 39301 35235 39359 35241
rect 41966 35232 41972 35284
rect 42024 35272 42030 35284
rect 47302 35272 47308 35284
rect 42024 35244 43024 35272
rect 47263 35244 47308 35272
rect 42024 35232 42030 35244
rect 38194 35204 38200 35216
rect 34287 35176 35848 35204
rect 37016 35176 38200 35204
rect 34287 35173 34299 35176
rect 34241 35167 34299 35173
rect 28813 35139 28871 35145
rect 28813 35105 28825 35139
rect 28859 35136 28871 35139
rect 28902 35136 28908 35148
rect 28859 35108 28908 35136
rect 28859 35105 28871 35108
rect 28813 35099 28871 35105
rect 28902 35096 28908 35108
rect 28960 35096 28966 35148
rect 33980 35136 34008 35164
rect 31220 35108 32628 35136
rect 28994 35068 29000 35080
rect 28955 35040 29000 35068
rect 28994 35028 29000 35040
rect 29052 35028 29058 35080
rect 30469 35071 30527 35077
rect 30469 35037 30481 35071
rect 30515 35037 30527 35071
rect 30650 35068 30656 35080
rect 30611 35040 30656 35068
rect 30469 35031 30527 35037
rect 27338 34960 27344 35012
rect 27396 35000 27402 35012
rect 27801 35003 27859 35009
rect 27801 35000 27813 35003
rect 27396 34972 27813 35000
rect 27396 34960 27402 34972
rect 27801 34969 27813 34972
rect 27847 35000 27859 35003
rect 30484 35000 30512 35031
rect 30650 35028 30656 35040
rect 30708 35028 30714 35080
rect 31220 35012 31248 35108
rect 31294 35028 31300 35080
rect 31352 35068 31358 35080
rect 31352 35040 31397 35068
rect 31352 35028 31358 35040
rect 31754 35028 31760 35080
rect 31812 35068 31818 35080
rect 32398 35068 32404 35080
rect 31812 35040 32404 35068
rect 31812 35028 31818 35040
rect 32398 35028 32404 35040
rect 32456 35028 32462 35080
rect 31202 35000 31208 35012
rect 27847 34972 28994 35000
rect 30484 34972 31208 35000
rect 27847 34969 27859 34972
rect 27801 34963 27859 34969
rect 28966 34932 28994 34972
rect 31202 34960 31208 34972
rect 31260 34960 31266 35012
rect 31849 35003 31907 35009
rect 31849 34969 31861 35003
rect 31895 35000 31907 35003
rect 32030 35000 32036 35012
rect 31895 34972 32036 35000
rect 31895 34969 31907 34972
rect 31849 34963 31907 34969
rect 32030 34960 32036 34972
rect 32088 34960 32094 35012
rect 32600 35000 32628 35108
rect 33428 35108 34008 35136
rect 34348 35108 36032 35136
rect 32766 35068 32772 35080
rect 32727 35040 32772 35068
rect 32766 35028 32772 35040
rect 32824 35028 32830 35080
rect 32953 35071 33011 35077
rect 32953 35037 32965 35071
rect 32999 35068 33011 35071
rect 33318 35068 33324 35080
rect 32999 35040 33324 35068
rect 32999 35037 33011 35040
rect 32953 35031 33011 35037
rect 32968 35000 32996 35031
rect 33318 35028 33324 35040
rect 33376 35028 33382 35080
rect 33428 35009 33456 35108
rect 33686 35068 33692 35080
rect 33647 35040 33692 35068
rect 33686 35028 33692 35040
rect 33744 35068 33750 35080
rect 34348 35068 34376 35108
rect 33744 35040 34376 35068
rect 35621 35071 35679 35077
rect 33744 35028 33750 35040
rect 35621 35037 35633 35071
rect 35667 35037 35679 35071
rect 35621 35031 35679 35037
rect 32600 34972 32996 35000
rect 33413 35003 33471 35009
rect 33413 34969 33425 35003
rect 33459 34969 33471 35003
rect 33413 34963 33471 34969
rect 33597 35003 33655 35009
rect 33597 34969 33609 35003
rect 33643 35000 33655 35003
rect 33778 35000 33784 35012
rect 33643 34972 33784 35000
rect 33643 34969 33655 34972
rect 33597 34963 33655 34969
rect 33778 34960 33784 34972
rect 33836 34960 33842 35012
rect 35636 35000 35664 35031
rect 35710 35028 35716 35080
rect 35768 35068 35774 35080
rect 35897 35071 35955 35077
rect 35897 35068 35909 35071
rect 35768 35040 35909 35068
rect 35768 35028 35774 35040
rect 35897 35037 35909 35040
rect 35943 35037 35955 35071
rect 36004 35068 36032 35108
rect 36170 35096 36176 35148
rect 36228 35136 36234 35148
rect 37016 35136 37044 35176
rect 38194 35164 38200 35176
rect 38252 35204 38258 35216
rect 38654 35204 38660 35216
rect 38252 35176 38660 35204
rect 38252 35164 38258 35176
rect 38654 35164 38660 35176
rect 38712 35164 38718 35216
rect 42996 35204 43024 35244
rect 47302 35232 47308 35244
rect 47360 35232 47366 35284
rect 49694 35272 49700 35284
rect 49655 35244 49700 35272
rect 49694 35232 49700 35244
rect 49752 35232 49758 35284
rect 52181 35275 52239 35281
rect 52181 35241 52193 35275
rect 52227 35272 52239 35275
rect 52546 35272 52552 35284
rect 52227 35244 52552 35272
rect 52227 35241 52239 35244
rect 52181 35235 52239 35241
rect 52546 35232 52552 35244
rect 52604 35272 52610 35284
rect 52733 35275 52791 35281
rect 52733 35272 52745 35275
rect 52604 35244 52745 35272
rect 52604 35232 52610 35244
rect 52733 35241 52745 35244
rect 52779 35241 52791 35275
rect 53650 35272 53656 35284
rect 53611 35244 53656 35272
rect 52733 35235 52791 35241
rect 53650 35232 53656 35244
rect 53708 35232 53714 35284
rect 42996 35176 43484 35204
rect 37182 35136 37188 35148
rect 36228 35108 37044 35136
rect 37143 35108 37188 35136
rect 36228 35096 36234 35108
rect 37016 35080 37044 35108
rect 37182 35096 37188 35108
rect 37240 35096 37246 35148
rect 37458 35136 37464 35148
rect 37292 35108 37464 35136
rect 36004 35040 36952 35068
rect 35897 35031 35955 35037
rect 36170 35000 36176 35012
rect 35636 34972 36176 35000
rect 36170 34960 36176 34972
rect 36228 34960 36234 35012
rect 36924 35000 36952 35040
rect 36998 35028 37004 35080
rect 37056 35068 37062 35080
rect 37292 35077 37320 35108
rect 37458 35096 37464 35108
rect 37516 35096 37522 35148
rect 38749 35139 38807 35145
rect 38749 35136 38761 35139
rect 37568 35108 38761 35136
rect 37568 35077 37596 35108
rect 38749 35105 38761 35108
rect 38795 35105 38807 35139
rect 38749 35099 38807 35105
rect 42705 35139 42763 35145
rect 42705 35105 42717 35139
rect 42751 35136 42763 35139
rect 43254 35136 43260 35148
rect 42751 35108 43260 35136
rect 42751 35105 42763 35108
rect 42705 35099 42763 35105
rect 43254 35096 43260 35108
rect 43312 35096 43318 35148
rect 43456 35136 43484 35176
rect 43530 35164 43536 35216
rect 43588 35204 43594 35216
rect 43717 35207 43775 35213
rect 43717 35204 43729 35207
rect 43588 35176 43729 35204
rect 43588 35164 43594 35176
rect 43717 35173 43729 35176
rect 43763 35173 43775 35207
rect 43717 35167 43775 35173
rect 49050 35164 49056 35216
rect 49108 35204 49114 35216
rect 49145 35207 49203 35213
rect 49145 35204 49157 35207
rect 49108 35176 49157 35204
rect 49108 35164 49114 35176
rect 49145 35173 49157 35176
rect 49191 35204 49203 35207
rect 53742 35204 53748 35216
rect 49191 35176 53748 35204
rect 49191 35173 49203 35176
rect 49145 35167 49203 35173
rect 43456 35108 45876 35136
rect 37277 35071 37335 35077
rect 37056 35040 37149 35068
rect 37056 35028 37062 35040
rect 37277 35037 37289 35071
rect 37323 35037 37335 35071
rect 37277 35031 37335 35037
rect 37369 35071 37427 35077
rect 37369 35037 37381 35071
rect 37415 35037 37427 35071
rect 37369 35031 37427 35037
rect 37553 35071 37611 35077
rect 37553 35037 37565 35071
rect 37599 35037 37611 35071
rect 37553 35031 37611 35037
rect 37292 35000 37320 35031
rect 36924 34972 37320 35000
rect 37384 35000 37412 35031
rect 37734 35028 37740 35080
rect 37792 35068 37798 35080
rect 38013 35071 38071 35077
rect 38013 35068 38025 35071
rect 37792 35040 38025 35068
rect 37792 35028 37798 35040
rect 38013 35037 38025 35040
rect 38059 35037 38071 35071
rect 38194 35068 38200 35080
rect 38155 35040 38200 35068
rect 38013 35031 38071 35037
rect 38194 35028 38200 35040
rect 38252 35028 38258 35080
rect 38657 35071 38715 35077
rect 38657 35037 38669 35071
rect 38703 35037 38715 35071
rect 38657 35031 38715 35037
rect 38841 35071 38899 35077
rect 38841 35037 38853 35071
rect 38887 35068 38899 35071
rect 38930 35068 38936 35080
rect 38887 35040 38936 35068
rect 38887 35037 38899 35040
rect 38841 35031 38899 35037
rect 37642 35000 37648 35012
rect 37384 34972 37648 35000
rect 37642 34960 37648 34972
rect 37700 35000 37706 35012
rect 38105 35003 38163 35009
rect 38105 35000 38117 35003
rect 37700 34972 38117 35000
rect 37700 34960 37706 34972
rect 38105 34969 38117 34972
rect 38151 34969 38163 35003
rect 38672 35000 38700 35031
rect 38930 35028 38936 35040
rect 38988 35028 38994 35080
rect 40773 35071 40831 35077
rect 40773 35037 40785 35071
rect 40819 35068 40831 35071
rect 41138 35068 41144 35080
rect 40819 35040 41144 35068
rect 40819 35037 40831 35040
rect 40773 35031 40831 35037
rect 41138 35028 41144 35040
rect 41196 35028 41202 35080
rect 41414 35028 41420 35080
rect 41472 35068 41478 35080
rect 41693 35071 41751 35077
rect 41693 35068 41705 35071
rect 41472 35040 41705 35068
rect 41472 35028 41478 35040
rect 41693 35037 41705 35040
rect 41739 35037 41751 35071
rect 41874 35068 41880 35080
rect 41835 35040 41880 35068
rect 41693 35031 41751 35037
rect 40126 35000 40132 35012
rect 38672 34972 38884 35000
rect 40039 34972 40132 35000
rect 38105 34963 38163 34969
rect 38856 34944 38884 34972
rect 40126 34960 40132 34972
rect 40184 35000 40190 35012
rect 41506 35000 41512 35012
rect 40184 34972 41512 35000
rect 40184 34960 40190 34972
rect 41506 34960 41512 34972
rect 41564 34960 41570 35012
rect 41708 35000 41736 35031
rect 41874 35028 41880 35040
rect 41932 35028 41938 35080
rect 42061 35071 42119 35077
rect 42061 35037 42073 35071
rect 42107 35068 42119 35071
rect 42797 35071 42855 35077
rect 42797 35068 42809 35071
rect 42107 35040 42809 35068
rect 42107 35037 42119 35040
rect 42061 35031 42119 35037
rect 42797 35037 42809 35040
rect 42843 35068 42855 35071
rect 43162 35068 43168 35080
rect 42843 35040 43168 35068
rect 42843 35037 42855 35040
rect 42797 35031 42855 35037
rect 43162 35028 43168 35040
rect 43220 35028 43226 35080
rect 43990 35068 43996 35080
rect 43951 35040 43996 35068
rect 43990 35028 43996 35040
rect 44048 35028 44054 35080
rect 42334 35000 42340 35012
rect 41708 34972 42340 35000
rect 42334 34960 42340 34972
rect 42392 35000 42398 35012
rect 42978 35000 42984 35012
rect 42392 34972 42984 35000
rect 42392 34960 42398 34972
rect 42978 34960 42984 34972
rect 43036 34960 43042 35012
rect 43717 35003 43775 35009
rect 43717 35000 43729 35003
rect 43272 34972 43729 35000
rect 30466 34932 30472 34944
rect 28966 34904 30472 34932
rect 30466 34892 30472 34904
rect 30524 34932 30530 34944
rect 32674 34932 32680 34944
rect 30524 34904 32680 34932
rect 30524 34892 30530 34904
rect 32674 34892 32680 34904
rect 32732 34892 32738 34944
rect 34514 34892 34520 34944
rect 34572 34932 34578 34944
rect 35434 34932 35440 34944
rect 34572 34904 35440 34932
rect 34572 34892 34578 34904
rect 35434 34892 35440 34904
rect 35492 34892 35498 34944
rect 35802 34932 35808 34944
rect 35763 34904 35808 34932
rect 35802 34892 35808 34904
rect 35860 34892 35866 34944
rect 36817 34935 36875 34941
rect 36817 34901 36829 34935
rect 36863 34932 36875 34935
rect 37550 34932 37556 34944
rect 36863 34904 37556 34932
rect 36863 34901 36875 34904
rect 36817 34895 36875 34901
rect 37550 34892 37556 34904
rect 37608 34892 37614 34944
rect 38838 34892 38844 34944
rect 38896 34892 38902 34944
rect 40957 34935 41015 34941
rect 40957 34901 40969 34935
rect 41003 34932 41015 34935
rect 41690 34932 41696 34944
rect 41003 34904 41696 34932
rect 41003 34901 41015 34904
rect 40957 34895 41015 34901
rect 41690 34892 41696 34904
rect 41748 34892 41754 34944
rect 42518 34892 42524 34944
rect 42576 34932 42582 34944
rect 43272 34941 43300 34972
rect 43717 34969 43729 34972
rect 43763 34969 43775 35003
rect 45848 35000 45876 35108
rect 45922 35096 45928 35148
rect 45980 35136 45986 35148
rect 47854 35136 47860 35148
rect 45980 35108 47860 35136
rect 45980 35096 45986 35108
rect 46658 35068 46664 35080
rect 46619 35040 46664 35068
rect 46658 35028 46664 35040
rect 46716 35028 46722 35080
rect 46768 35077 46796 35108
rect 47854 35096 47860 35108
rect 47912 35136 47918 35148
rect 47912 35108 48268 35136
rect 47912 35096 47918 35108
rect 46754 35071 46812 35077
rect 46754 35037 46766 35071
rect 46800 35037 46812 35071
rect 46934 35068 46940 35080
rect 46895 35040 46940 35068
rect 46754 35031 46812 35037
rect 46934 35028 46940 35040
rect 46992 35028 46998 35080
rect 47167 35071 47225 35077
rect 47167 35037 47179 35071
rect 47213 35068 47225 35071
rect 48130 35068 48136 35080
rect 47213 35040 48136 35068
rect 47213 35037 47225 35040
rect 47167 35031 47225 35037
rect 48130 35028 48136 35040
rect 48188 35028 48194 35080
rect 48240 35068 48268 35108
rect 48314 35096 48320 35148
rect 48372 35136 48378 35148
rect 53576 35145 53604 35176
rect 53742 35164 53748 35176
rect 53800 35164 53806 35216
rect 55766 35164 55772 35216
rect 55824 35204 55830 35216
rect 56594 35204 56600 35216
rect 55824 35176 56600 35204
rect 55824 35164 55830 35176
rect 56594 35164 56600 35176
rect 56652 35204 56658 35216
rect 57885 35207 57943 35213
rect 57885 35204 57897 35207
rect 56652 35176 57897 35204
rect 56652 35164 56658 35176
rect 57885 35173 57897 35176
rect 57931 35204 57943 35207
rect 58066 35204 58072 35216
rect 57931 35176 58072 35204
rect 57931 35173 57943 35176
rect 57885 35167 57943 35173
rect 58066 35164 58072 35176
rect 58124 35164 58130 35216
rect 50525 35139 50583 35145
rect 50525 35136 50537 35139
rect 48372 35108 50537 35136
rect 48372 35096 48378 35108
rect 50525 35105 50537 35108
rect 50571 35105 50583 35139
rect 50525 35099 50583 35105
rect 53561 35139 53619 35145
rect 53561 35105 53573 35139
rect 53607 35105 53619 35139
rect 54849 35139 54907 35145
rect 54849 35136 54861 35139
rect 53561 35099 53619 35105
rect 53668 35108 54861 35136
rect 48593 35071 48651 35077
rect 48593 35068 48605 35071
rect 48240 35040 48605 35068
rect 48593 35037 48605 35040
rect 48639 35068 48651 35071
rect 48682 35068 48688 35080
rect 48639 35040 48688 35068
rect 48639 35037 48651 35040
rect 48593 35031 48651 35037
rect 48682 35028 48688 35040
rect 48740 35028 48746 35080
rect 48866 35068 48872 35080
rect 48827 35040 48872 35068
rect 48866 35028 48872 35040
rect 48924 35028 48930 35080
rect 49237 35071 49295 35077
rect 49237 35037 49249 35071
rect 49283 35037 49295 35071
rect 50798 35068 50804 35080
rect 50759 35040 50804 35068
rect 49237 35031 49295 35037
rect 47029 35003 47087 35009
rect 47029 35000 47041 35003
rect 45848 34972 47041 35000
rect 43717 34963 43775 34969
rect 47029 34969 47041 34972
rect 47075 35000 47087 35003
rect 47578 35000 47584 35012
rect 47075 34972 47584 35000
rect 47075 34969 47087 34972
rect 47029 34963 47087 34969
rect 47578 34960 47584 34972
rect 47636 34960 47642 35012
rect 48314 34960 48320 35012
rect 48372 35000 48378 35012
rect 48774 35000 48780 35012
rect 48372 34972 48780 35000
rect 48372 34960 48378 34972
rect 48774 34960 48780 34972
rect 48832 35000 48838 35012
rect 49252 35000 49280 35031
rect 50798 35028 50804 35040
rect 50856 35028 50862 35080
rect 53190 35028 53196 35080
rect 53248 35068 53254 35080
rect 53668 35068 53696 35108
rect 54849 35105 54861 35108
rect 54895 35105 54907 35139
rect 54849 35099 54907 35105
rect 53248 35040 53696 35068
rect 53745 35071 53803 35077
rect 53248 35028 53254 35040
rect 53745 35037 53757 35071
rect 53791 35037 53803 35071
rect 53745 35031 53803 35037
rect 53837 35071 53895 35077
rect 53837 35037 53849 35071
rect 53883 35068 53895 35071
rect 54754 35068 54760 35080
rect 53883 35040 54760 35068
rect 53883 35037 53895 35040
rect 53837 35031 53895 35037
rect 48832 34972 49280 35000
rect 48832 34960 48838 34972
rect 49970 34960 49976 35012
rect 50028 35000 50034 35012
rect 53374 35000 53380 35012
rect 50028 34972 53380 35000
rect 50028 34960 50034 34972
rect 53374 34960 53380 34972
rect 53432 35000 53438 35012
rect 53760 35000 53788 35031
rect 54754 35028 54760 35040
rect 54812 35028 54818 35080
rect 53432 34972 53788 35000
rect 54864 35000 54892 35099
rect 55490 35096 55496 35148
rect 55548 35136 55554 35148
rect 57425 35139 57483 35145
rect 57425 35136 57437 35139
rect 55548 35108 57437 35136
rect 55548 35096 55554 35108
rect 57425 35105 57437 35108
rect 57471 35136 57483 35139
rect 57974 35136 57980 35148
rect 57471 35108 57980 35136
rect 57471 35105 57483 35108
rect 57425 35099 57483 35105
rect 57974 35096 57980 35108
rect 58032 35096 58038 35148
rect 55766 35028 55772 35080
rect 55824 35068 55830 35080
rect 55953 35071 56011 35077
rect 55953 35068 55965 35071
rect 55824 35040 55965 35068
rect 55824 35028 55830 35040
rect 55953 35037 55965 35040
rect 55999 35037 56011 35071
rect 56134 35068 56140 35080
rect 56095 35040 56140 35068
rect 55953 35031 56011 35037
rect 56134 35028 56140 35040
rect 56192 35028 56198 35080
rect 56229 35071 56287 35077
rect 56229 35037 56241 35071
rect 56275 35068 56287 35071
rect 56318 35068 56324 35080
rect 56275 35040 56324 35068
rect 56275 35037 56287 35040
rect 56229 35031 56287 35037
rect 56318 35028 56324 35040
rect 56376 35028 56382 35080
rect 57146 35068 57152 35080
rect 57107 35040 57152 35068
rect 57146 35028 57152 35040
rect 57204 35028 57210 35080
rect 57330 35068 57336 35080
rect 57291 35040 57336 35068
rect 57330 35028 57336 35040
rect 57388 35028 57394 35080
rect 57698 35000 57704 35012
rect 54864 34972 57704 35000
rect 53432 34960 53438 34972
rect 57698 34960 57704 34972
rect 57756 34960 57762 35012
rect 42889 34935 42947 34941
rect 42889 34932 42901 34935
rect 42576 34904 42901 34932
rect 42576 34892 42582 34904
rect 42889 34901 42901 34904
rect 42935 34901 42947 34935
rect 42889 34895 42947 34901
rect 43257 34935 43315 34941
rect 43257 34901 43269 34935
rect 43303 34901 43315 34935
rect 43898 34932 43904 34944
rect 43859 34904 43904 34932
rect 43257 34895 43315 34901
rect 43898 34892 43904 34904
rect 43956 34892 43962 34944
rect 44450 34932 44456 34944
rect 44411 34904 44456 34932
rect 44450 34892 44456 34904
rect 44508 34892 44514 34944
rect 45186 34892 45192 34944
rect 45244 34932 45250 34944
rect 45281 34935 45339 34941
rect 45281 34932 45293 34935
rect 45244 34904 45293 34932
rect 45244 34892 45250 34904
rect 45281 34901 45293 34904
rect 45327 34932 45339 34935
rect 46934 34932 46940 34944
rect 45327 34904 46940 34932
rect 45327 34901 45339 34904
rect 45281 34895 45339 34901
rect 46934 34892 46940 34904
rect 46992 34892 46998 34944
rect 47857 34935 47915 34941
rect 47857 34901 47869 34935
rect 47903 34932 47915 34935
rect 47946 34932 47952 34944
rect 47903 34904 47952 34932
rect 47903 34901 47915 34904
rect 47857 34895 47915 34901
rect 47946 34892 47952 34904
rect 48004 34892 48010 34944
rect 51350 34892 51356 34944
rect 51408 34932 51414 34944
rect 51445 34935 51503 34941
rect 51445 34932 51457 34935
rect 51408 34904 51457 34932
rect 51408 34892 51414 34904
rect 51445 34901 51457 34904
rect 51491 34901 51503 34935
rect 51445 34895 51503 34901
rect 52638 34892 52644 34944
rect 52696 34932 52702 34944
rect 54110 34932 54116 34944
rect 52696 34904 54116 34932
rect 52696 34892 52702 34904
rect 54110 34892 54116 34904
rect 54168 34932 54174 34944
rect 54297 34935 54355 34941
rect 54297 34932 54309 34935
rect 54168 34904 54309 34932
rect 54168 34892 54174 34904
rect 54297 34901 54309 34904
rect 54343 34901 54355 34935
rect 54297 34895 54355 34901
rect 55769 34935 55827 34941
rect 55769 34901 55781 34935
rect 55815 34932 55827 34935
rect 55950 34932 55956 34944
rect 55815 34904 55956 34932
rect 55815 34901 55827 34904
rect 55769 34895 55827 34901
rect 55950 34892 55956 34904
rect 56008 34892 56014 34944
rect 56962 34932 56968 34944
rect 56923 34904 56968 34932
rect 56962 34892 56968 34904
rect 57020 34892 57026 34944
rect 1104 34842 58880 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 58880 34842
rect 1104 34768 58880 34790
rect 27525 34731 27583 34737
rect 27525 34697 27537 34731
rect 27571 34728 27583 34731
rect 27614 34728 27620 34740
rect 27571 34700 27620 34728
rect 27571 34697 27583 34700
rect 27525 34691 27583 34697
rect 27614 34688 27620 34700
rect 27672 34688 27678 34740
rect 28994 34688 29000 34740
rect 29052 34728 29058 34740
rect 32490 34728 32496 34740
rect 29052 34700 31892 34728
rect 32451 34700 32496 34728
rect 29052 34688 29058 34700
rect 29086 34620 29092 34672
rect 29144 34620 29150 34672
rect 30101 34663 30159 34669
rect 30101 34629 30113 34663
rect 30147 34660 30159 34663
rect 30190 34660 30196 34672
rect 30147 34632 30196 34660
rect 30147 34629 30159 34632
rect 30101 34623 30159 34629
rect 30190 34620 30196 34632
rect 30248 34620 30254 34672
rect 30650 34620 30656 34672
rect 30708 34660 30714 34672
rect 31754 34660 31760 34672
rect 30708 34632 31340 34660
rect 30708 34620 30714 34632
rect 27338 34592 27344 34604
rect 27299 34564 27344 34592
rect 27338 34552 27344 34564
rect 27396 34552 27402 34604
rect 31113 34595 31171 34601
rect 31113 34561 31125 34595
rect 31159 34592 31171 34595
rect 31202 34592 31208 34604
rect 31159 34564 31208 34592
rect 31159 34561 31171 34564
rect 31113 34555 31171 34561
rect 31202 34552 31208 34564
rect 31260 34552 31266 34604
rect 31312 34601 31340 34632
rect 31726 34620 31760 34660
rect 31812 34620 31818 34672
rect 31297 34595 31355 34601
rect 31297 34561 31309 34595
rect 31343 34561 31355 34595
rect 31297 34555 31355 34561
rect 31573 34595 31631 34601
rect 31573 34561 31585 34595
rect 31619 34592 31631 34595
rect 31726 34592 31754 34620
rect 31619 34564 31754 34592
rect 31619 34561 31631 34564
rect 31573 34555 31631 34561
rect 28074 34524 28080 34536
rect 28035 34496 28080 34524
rect 28074 34484 28080 34496
rect 28132 34484 28138 34536
rect 31312 34524 31340 34555
rect 31662 34524 31668 34536
rect 31312 34496 31668 34524
rect 31662 34484 31668 34496
rect 31720 34484 31726 34536
rect 31757 34527 31815 34533
rect 31757 34493 31769 34527
rect 31803 34524 31815 34527
rect 31864 34524 31892 34700
rect 32490 34688 32496 34700
rect 32548 34688 32554 34740
rect 32674 34688 32680 34740
rect 32732 34728 32738 34740
rect 32732 34700 40908 34728
rect 32732 34688 32738 34700
rect 31938 34620 31944 34672
rect 31996 34660 32002 34672
rect 33226 34660 33232 34672
rect 31996 34632 33232 34660
rect 31996 34620 32002 34632
rect 32324 34601 32352 34632
rect 33226 34620 33232 34632
rect 33284 34620 33290 34672
rect 35253 34663 35311 34669
rect 35253 34629 35265 34663
rect 35299 34660 35311 34663
rect 35342 34660 35348 34672
rect 35299 34632 35348 34660
rect 35299 34629 35311 34632
rect 35253 34623 35311 34629
rect 35342 34620 35348 34632
rect 35400 34620 35406 34672
rect 36817 34663 36875 34669
rect 36817 34629 36829 34663
rect 36863 34660 36875 34663
rect 36998 34660 37004 34672
rect 36863 34632 37004 34660
rect 36863 34629 36875 34632
rect 36817 34623 36875 34629
rect 36998 34620 37004 34632
rect 37056 34620 37062 34672
rect 38654 34660 38660 34672
rect 37384 34632 38660 34660
rect 32309 34595 32367 34601
rect 32309 34561 32321 34595
rect 32355 34561 32367 34595
rect 33134 34592 33140 34604
rect 33095 34564 33140 34592
rect 32309 34555 32367 34561
rect 33134 34552 33140 34564
rect 33192 34552 33198 34604
rect 33778 34592 33784 34604
rect 33739 34564 33784 34592
rect 33778 34552 33784 34564
rect 33836 34592 33842 34604
rect 34793 34595 34851 34601
rect 34793 34592 34805 34595
rect 33836 34564 34805 34592
rect 33836 34552 33842 34564
rect 34793 34561 34805 34564
rect 34839 34561 34851 34595
rect 34793 34555 34851 34561
rect 35437 34595 35495 34601
rect 35437 34561 35449 34595
rect 35483 34561 35495 34595
rect 35437 34555 35495 34561
rect 33873 34527 33931 34533
rect 33873 34524 33885 34527
rect 31803 34496 33885 34524
rect 31803 34493 31815 34496
rect 31757 34487 31815 34493
rect 33873 34493 33885 34496
rect 33919 34493 33931 34527
rect 33873 34487 33931 34493
rect 34330 34484 34336 34536
rect 34388 34524 34394 34536
rect 34701 34527 34759 34533
rect 34701 34524 34713 34527
rect 34388 34496 34713 34524
rect 34388 34484 34394 34496
rect 34701 34493 34713 34496
rect 34747 34493 34759 34527
rect 34701 34487 34759 34493
rect 35342 34484 35348 34536
rect 35400 34524 35406 34536
rect 35452 34524 35480 34555
rect 35526 34552 35532 34604
rect 35584 34592 35590 34604
rect 36265 34595 36323 34601
rect 35584 34564 35629 34592
rect 35584 34552 35590 34564
rect 36265 34561 36277 34595
rect 36311 34592 36323 34595
rect 37384 34592 37412 34632
rect 38654 34620 38660 34632
rect 38712 34620 38718 34672
rect 39298 34620 39304 34672
rect 39356 34620 39362 34672
rect 40310 34660 40316 34672
rect 40271 34632 40316 34660
rect 40310 34620 40316 34632
rect 40368 34620 40374 34672
rect 40880 34669 40908 34700
rect 41046 34688 41052 34740
rect 41104 34728 41110 34740
rect 42334 34728 42340 34740
rect 41104 34700 42340 34728
rect 41104 34688 41110 34700
rect 42334 34688 42340 34700
rect 42392 34728 42398 34740
rect 42613 34731 42671 34737
rect 42613 34728 42625 34731
rect 42392 34700 42625 34728
rect 42392 34688 42398 34700
rect 42613 34697 42625 34700
rect 42659 34728 42671 34731
rect 43714 34728 43720 34740
rect 42659 34700 43720 34728
rect 42659 34697 42671 34700
rect 42613 34691 42671 34697
rect 43714 34688 43720 34700
rect 43772 34728 43778 34740
rect 44450 34728 44456 34740
rect 43772 34700 44456 34728
rect 43772 34688 43778 34700
rect 44450 34688 44456 34700
rect 44508 34688 44514 34740
rect 48777 34731 48835 34737
rect 48777 34697 48789 34731
rect 48823 34728 48835 34731
rect 48958 34728 48964 34740
rect 48823 34700 48964 34728
rect 48823 34697 48835 34700
rect 48777 34691 48835 34697
rect 48958 34688 48964 34700
rect 49016 34728 49022 34740
rect 50982 34728 50988 34740
rect 49016 34700 50988 34728
rect 49016 34688 49022 34700
rect 50982 34688 50988 34700
rect 51040 34688 51046 34740
rect 56318 34728 56324 34740
rect 54036 34700 56324 34728
rect 40865 34663 40923 34669
rect 40865 34629 40877 34663
rect 40911 34660 40923 34663
rect 44269 34663 44327 34669
rect 44269 34660 44281 34663
rect 40911 34632 44281 34660
rect 40911 34629 40923 34632
rect 40865 34623 40923 34629
rect 44269 34629 44281 34632
rect 44315 34629 44327 34663
rect 45922 34660 45928 34672
rect 44269 34623 44327 34629
rect 45020 34632 45928 34660
rect 36311 34564 37412 34592
rect 37461 34595 37519 34601
rect 36311 34561 36323 34564
rect 36265 34555 36323 34561
rect 37461 34561 37473 34595
rect 37507 34561 37519 34595
rect 37461 34555 37519 34561
rect 37553 34595 37611 34601
rect 37553 34561 37565 34595
rect 37599 34592 37611 34595
rect 37642 34592 37648 34604
rect 37599 34564 37648 34592
rect 37599 34561 37611 34564
rect 37553 34555 37611 34561
rect 37182 34524 37188 34536
rect 35400 34496 35480 34524
rect 35544 34496 37188 34524
rect 35400 34484 35406 34496
rect 33321 34459 33379 34465
rect 33321 34425 33333 34459
rect 33367 34456 33379 34459
rect 33410 34456 33416 34468
rect 33367 34428 33416 34456
rect 33367 34425 33379 34428
rect 33321 34419 33379 34425
rect 33410 34416 33416 34428
rect 33468 34416 33474 34468
rect 28340 34391 28398 34397
rect 28340 34357 28352 34391
rect 28386 34388 28398 34391
rect 28534 34388 28540 34400
rect 28386 34360 28540 34388
rect 28386 34357 28398 34360
rect 28340 34351 28398 34357
rect 28534 34348 28540 34360
rect 28592 34348 28598 34400
rect 32306 34348 32312 34400
rect 32364 34388 32370 34400
rect 32766 34388 32772 34400
rect 32364 34360 32772 34388
rect 32364 34348 32370 34360
rect 32766 34348 32772 34360
rect 32824 34388 32830 34400
rect 33042 34388 33048 34400
rect 32824 34360 33048 34388
rect 32824 34348 32830 34360
rect 33042 34348 33048 34360
rect 33100 34388 33106 34400
rect 35544 34388 35572 34496
rect 37182 34484 37188 34496
rect 37240 34524 37246 34536
rect 37476 34524 37504 34555
rect 37642 34552 37648 34564
rect 37700 34552 37706 34604
rect 38286 34592 38292 34604
rect 38247 34564 38292 34592
rect 38286 34552 38292 34564
rect 38344 34552 38350 34604
rect 41693 34595 41751 34601
rect 41693 34561 41705 34595
rect 41739 34592 41751 34595
rect 41966 34592 41972 34604
rect 41739 34564 41972 34592
rect 41739 34561 41751 34564
rect 41693 34555 41751 34561
rect 41966 34552 41972 34564
rect 42024 34552 42030 34604
rect 43162 34552 43168 34604
rect 43220 34592 43226 34604
rect 43441 34595 43499 34601
rect 43441 34592 43453 34595
rect 43220 34564 43453 34592
rect 43220 34552 43226 34564
rect 43441 34561 43453 34564
rect 43487 34592 43499 34595
rect 44082 34592 44088 34604
rect 43487 34564 44088 34592
rect 43487 34561 43499 34564
rect 43441 34555 43499 34561
rect 44082 34552 44088 34564
rect 44140 34552 44146 34604
rect 45020 34601 45048 34632
rect 45922 34620 45928 34632
rect 45980 34620 45986 34672
rect 48866 34660 48872 34672
rect 47136 34632 48872 34660
rect 45005 34595 45063 34601
rect 45005 34561 45017 34595
rect 45051 34561 45063 34595
rect 45005 34555 45063 34561
rect 45830 34552 45836 34604
rect 45888 34592 45894 34604
rect 46017 34595 46075 34601
rect 46017 34592 46029 34595
rect 45888 34564 46029 34592
rect 45888 34552 45894 34564
rect 46017 34561 46029 34564
rect 46063 34561 46075 34595
rect 46017 34555 46075 34561
rect 46106 34552 46112 34604
rect 46164 34592 46170 34604
rect 46566 34592 46572 34604
rect 46164 34564 46572 34592
rect 46164 34552 46170 34564
rect 46566 34552 46572 34564
rect 46624 34592 46630 34604
rect 47029 34595 47087 34601
rect 47029 34592 47041 34595
rect 46624 34564 47041 34592
rect 46624 34552 46630 34564
rect 47029 34561 47041 34564
rect 47075 34561 47087 34595
rect 47029 34555 47087 34561
rect 37240 34496 37504 34524
rect 37737 34527 37795 34533
rect 37240 34484 37246 34496
rect 37737 34493 37749 34527
rect 37783 34524 37795 34527
rect 37826 34524 37832 34536
rect 37783 34496 37832 34524
rect 37783 34493 37795 34496
rect 37737 34487 37795 34493
rect 37826 34484 37832 34496
rect 37884 34484 37890 34536
rect 41046 34524 41052 34536
rect 41007 34496 41052 34524
rect 41046 34484 41052 34496
rect 41104 34484 41110 34536
rect 41138 34484 41144 34536
rect 41196 34524 41202 34536
rect 43530 34524 43536 34536
rect 41196 34496 41552 34524
rect 43491 34496 43536 34524
rect 41196 34484 41202 34496
rect 41524 34465 41552 34496
rect 43530 34484 43536 34496
rect 43588 34484 43594 34536
rect 45094 34524 45100 34536
rect 45055 34496 45100 34524
rect 45094 34484 45100 34496
rect 45152 34484 45158 34536
rect 45925 34527 45983 34533
rect 45925 34493 45937 34527
rect 45971 34493 45983 34527
rect 46845 34527 46903 34533
rect 46845 34524 46857 34527
rect 45925 34487 45983 34493
rect 46124 34496 46857 34524
rect 41509 34459 41567 34465
rect 41509 34425 41521 34459
rect 41555 34425 41567 34459
rect 41509 34419 41567 34425
rect 45373 34459 45431 34465
rect 45373 34425 45385 34459
rect 45419 34456 45431 34459
rect 45940 34456 45968 34487
rect 45419 34428 45968 34456
rect 45419 34425 45431 34428
rect 45373 34419 45431 34425
rect 36170 34388 36176 34400
rect 33100 34360 35572 34388
rect 36131 34360 36176 34388
rect 33100 34348 33106 34360
rect 36170 34348 36176 34360
rect 36228 34348 36234 34400
rect 37642 34348 37648 34400
rect 37700 34388 37706 34400
rect 38552 34391 38610 34397
rect 37700 34360 37745 34388
rect 37700 34348 37706 34360
rect 38552 34357 38564 34391
rect 38598 34388 38610 34391
rect 39114 34388 39120 34400
rect 38598 34360 39120 34388
rect 38598 34357 38610 34360
rect 38552 34351 38610 34357
rect 39114 34348 39120 34360
rect 39172 34348 39178 34400
rect 43717 34391 43775 34397
rect 43717 34357 43729 34391
rect 43763 34388 43775 34391
rect 44174 34388 44180 34400
rect 43763 34360 44180 34388
rect 43763 34357 43775 34360
rect 43717 34351 43775 34357
rect 44174 34348 44180 34360
rect 44232 34348 44238 34400
rect 44542 34348 44548 34400
rect 44600 34388 44606 34400
rect 46124 34388 46152 34496
rect 46845 34493 46857 34496
rect 46891 34524 46903 34527
rect 47136 34524 47164 34632
rect 48866 34620 48872 34632
rect 48924 34660 48930 34672
rect 49602 34660 49608 34672
rect 48924 34632 49608 34660
rect 48924 34620 48930 34632
rect 49602 34620 49608 34632
rect 49660 34620 49666 34672
rect 52362 34620 52368 34672
rect 52420 34660 52426 34672
rect 53101 34663 53159 34669
rect 53101 34660 53113 34663
rect 52420 34632 53113 34660
rect 52420 34620 52426 34632
rect 53101 34629 53113 34632
rect 53147 34629 53159 34663
rect 53101 34623 53159 34629
rect 47854 34552 47860 34604
rect 47912 34592 47918 34604
rect 47949 34595 48007 34601
rect 47949 34592 47961 34595
rect 47912 34564 47961 34592
rect 47912 34552 47918 34564
rect 47949 34561 47961 34564
rect 47995 34561 48007 34595
rect 47949 34555 48007 34561
rect 48314 34552 48320 34604
rect 48372 34592 48378 34604
rect 48501 34595 48559 34601
rect 48501 34592 48513 34595
rect 48372 34564 48513 34592
rect 48372 34552 48378 34564
rect 48501 34561 48513 34564
rect 48547 34561 48559 34595
rect 48501 34555 48559 34561
rect 48682 34552 48688 34604
rect 48740 34592 48746 34604
rect 48961 34595 49019 34601
rect 48961 34592 48973 34595
rect 48740 34564 48973 34592
rect 48740 34552 48746 34564
rect 48961 34561 48973 34564
rect 49007 34561 49019 34595
rect 49326 34592 49332 34604
rect 49287 34564 49332 34592
rect 48961 34555 49019 34561
rect 49326 34552 49332 34564
rect 49384 34552 49390 34604
rect 50798 34552 50804 34604
rect 50856 34592 50862 34604
rect 50985 34595 51043 34601
rect 50985 34592 50997 34595
rect 50856 34564 50997 34592
rect 50856 34552 50862 34564
rect 50985 34561 50997 34564
rect 51031 34561 51043 34595
rect 50985 34555 51043 34561
rect 51442 34552 51448 34604
rect 51500 34592 51506 34604
rect 51718 34592 51724 34604
rect 51500 34564 51724 34592
rect 51500 34552 51506 34564
rect 51718 34552 51724 34564
rect 51776 34552 51782 34604
rect 52914 34592 52920 34604
rect 52875 34564 52920 34592
rect 52914 34552 52920 34564
rect 52972 34552 52978 34604
rect 54036 34601 54064 34700
rect 56318 34688 56324 34700
rect 56376 34688 56382 34740
rect 57146 34688 57152 34740
rect 57204 34728 57210 34740
rect 58167 34731 58225 34737
rect 58167 34728 58179 34731
rect 57204 34700 58179 34728
rect 57204 34688 57210 34700
rect 58167 34697 58179 34700
rect 58213 34697 58225 34731
rect 58167 34691 58225 34697
rect 54570 34620 54576 34672
rect 54628 34660 54634 34672
rect 54628 34632 57192 34660
rect 54628 34620 54634 34632
rect 54021 34595 54079 34601
rect 54021 34561 54033 34595
rect 54067 34561 54079 34595
rect 55490 34592 55496 34604
rect 55451 34564 55496 34592
rect 54021 34555 54079 34561
rect 55490 34552 55496 34564
rect 55548 34552 55554 34604
rect 56318 34592 56324 34604
rect 56279 34564 56324 34592
rect 56318 34552 56324 34564
rect 56376 34552 56382 34604
rect 57164 34601 57192 34632
rect 57974 34620 57980 34672
rect 58032 34660 58038 34672
rect 58253 34663 58311 34669
rect 58253 34660 58265 34663
rect 58032 34632 58265 34660
rect 58032 34620 58038 34632
rect 58253 34629 58265 34632
rect 58299 34629 58311 34663
rect 58253 34623 58311 34629
rect 56505 34595 56563 34601
rect 56505 34561 56517 34595
rect 56551 34561 56563 34595
rect 56505 34555 56563 34561
rect 57149 34595 57207 34601
rect 57149 34561 57161 34595
rect 57195 34561 57207 34595
rect 58066 34592 58072 34604
rect 58027 34564 58072 34592
rect 57149 34555 57207 34561
rect 46891 34496 47164 34524
rect 47213 34527 47271 34533
rect 46891 34493 46903 34496
rect 46845 34487 46903 34493
rect 47213 34493 47225 34527
rect 47259 34524 47271 34527
rect 48700 34524 48728 34552
rect 47259 34496 48728 34524
rect 47259 34493 47271 34496
rect 47213 34487 47271 34493
rect 51534 34484 51540 34536
rect 51592 34524 51598 34536
rect 51629 34527 51687 34533
rect 51629 34524 51641 34527
rect 51592 34496 51641 34524
rect 51592 34484 51598 34496
rect 51629 34493 51641 34496
rect 51675 34524 51687 34527
rect 53929 34527 53987 34533
rect 53929 34524 53941 34527
rect 51675 34496 53941 34524
rect 51675 34493 51687 34496
rect 51629 34487 51687 34493
rect 53929 34493 53941 34496
rect 53975 34493 53987 34527
rect 55582 34524 55588 34536
rect 55543 34496 55588 34524
rect 53929 34487 53987 34493
rect 55582 34484 55588 34496
rect 55640 34484 55646 34536
rect 55861 34527 55919 34533
rect 55861 34493 55873 34527
rect 55907 34524 55919 34527
rect 56134 34524 56140 34536
rect 55907 34496 56140 34524
rect 55907 34493 55919 34496
rect 55861 34487 55919 34493
rect 56134 34484 56140 34496
rect 56192 34524 56198 34536
rect 56520 34524 56548 34555
rect 58066 34552 58072 34564
rect 58124 34552 58130 34604
rect 58345 34595 58403 34601
rect 58345 34561 58357 34595
rect 58391 34561 58403 34595
rect 58345 34555 58403 34561
rect 57054 34524 57060 34536
rect 56192 34496 56548 34524
rect 57015 34496 57060 34524
rect 56192 34484 56198 34496
rect 57054 34484 57060 34496
rect 57112 34484 57118 34536
rect 58360 34524 58388 34555
rect 57440 34496 58388 34524
rect 52089 34459 52147 34465
rect 52089 34425 52101 34459
rect 52135 34456 52147 34459
rect 52454 34456 52460 34468
rect 52135 34428 52460 34456
rect 52135 34425 52147 34428
rect 52089 34419 52147 34425
rect 52454 34416 52460 34428
rect 52512 34456 52518 34468
rect 52914 34456 52920 34468
rect 52512 34428 52920 34456
rect 52512 34416 52518 34428
rect 52914 34416 52920 34428
rect 52972 34416 52978 34468
rect 46290 34388 46296 34400
rect 44600 34360 46152 34388
rect 46251 34360 46296 34388
rect 44600 34348 44606 34360
rect 46290 34348 46296 34360
rect 46348 34348 46354 34400
rect 47854 34388 47860 34400
rect 47815 34360 47860 34388
rect 47854 34348 47860 34360
rect 47912 34348 47918 34400
rect 49970 34348 49976 34400
rect 50028 34388 50034 34400
rect 50433 34391 50491 34397
rect 50433 34388 50445 34391
rect 50028 34360 50445 34388
rect 50028 34348 50034 34360
rect 50433 34357 50445 34360
rect 50479 34357 50491 34391
rect 50433 34351 50491 34357
rect 53285 34391 53343 34397
rect 53285 34357 53297 34391
rect 53331 34388 53343 34391
rect 53374 34388 53380 34400
rect 53331 34360 53380 34388
rect 53331 34357 53343 34360
rect 53285 34351 53343 34357
rect 53374 34348 53380 34360
rect 53432 34348 53438 34400
rect 54389 34391 54447 34397
rect 54389 34357 54401 34391
rect 54435 34388 54447 34391
rect 54478 34388 54484 34400
rect 54435 34360 54484 34388
rect 54435 34357 54447 34360
rect 54389 34351 54447 34357
rect 54478 34348 54484 34360
rect 54536 34348 54542 34400
rect 56042 34348 56048 34400
rect 56100 34388 56106 34400
rect 56413 34391 56471 34397
rect 56413 34388 56425 34391
rect 56100 34360 56425 34388
rect 56100 34348 56106 34360
rect 56413 34357 56425 34360
rect 56459 34357 56471 34391
rect 56413 34351 56471 34357
rect 57330 34348 57336 34400
rect 57388 34388 57394 34400
rect 57440 34397 57468 34496
rect 57425 34391 57483 34397
rect 57425 34388 57437 34391
rect 57388 34360 57437 34388
rect 57388 34348 57394 34360
rect 57425 34357 57437 34360
rect 57471 34357 57483 34391
rect 57425 34351 57483 34357
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 28074 34144 28080 34196
rect 28132 34184 28138 34196
rect 28261 34187 28319 34193
rect 28261 34184 28273 34187
rect 28132 34156 28273 34184
rect 28132 34144 28138 34156
rect 28261 34153 28273 34156
rect 28307 34153 28319 34187
rect 29086 34184 29092 34196
rect 29047 34156 29092 34184
rect 28261 34147 28319 34153
rect 29086 34144 29092 34156
rect 29144 34144 29150 34196
rect 29733 34187 29791 34193
rect 29733 34153 29745 34187
rect 29779 34184 29791 34187
rect 30650 34184 30656 34196
rect 29779 34156 30656 34184
rect 29779 34153 29791 34156
rect 29733 34147 29791 34153
rect 30650 34144 30656 34156
rect 30708 34144 30714 34196
rect 31223 34187 31281 34193
rect 31223 34153 31235 34187
rect 31269 34184 31281 34187
rect 33045 34187 33103 34193
rect 31269 34156 31754 34184
rect 31269 34153 31281 34156
rect 31223 34147 31281 34153
rect 31726 34116 31754 34156
rect 33045 34153 33057 34187
rect 33091 34184 33103 34187
rect 33134 34184 33140 34196
rect 33091 34156 33140 34184
rect 33091 34153 33103 34156
rect 33045 34147 33103 34153
rect 33134 34144 33140 34156
rect 33192 34144 33198 34196
rect 36354 34184 36360 34196
rect 33336 34156 36360 34184
rect 33336 34116 33364 34156
rect 36354 34144 36360 34156
rect 36412 34144 36418 34196
rect 36633 34187 36691 34193
rect 36633 34153 36645 34187
rect 36679 34184 36691 34187
rect 37366 34184 37372 34196
rect 36679 34156 37372 34184
rect 36679 34153 36691 34156
rect 36633 34147 36691 34153
rect 37366 34144 37372 34156
rect 37424 34144 37430 34196
rect 39298 34144 39304 34196
rect 39356 34184 39362 34196
rect 39393 34187 39451 34193
rect 39393 34184 39405 34187
rect 39356 34156 39405 34184
rect 39356 34144 39362 34156
rect 39393 34153 39405 34156
rect 39439 34153 39451 34187
rect 43254 34184 43260 34196
rect 43215 34156 43260 34184
rect 39393 34147 39451 34153
rect 43254 34144 43260 34156
rect 43312 34144 43318 34196
rect 43898 34144 43904 34196
rect 43956 34184 43962 34196
rect 45830 34184 45836 34196
rect 43956 34156 45836 34184
rect 43956 34144 43962 34156
rect 45830 34144 45836 34156
rect 45888 34184 45894 34196
rect 48590 34184 48596 34196
rect 45888 34156 48596 34184
rect 45888 34144 45894 34156
rect 48590 34144 48596 34156
rect 48648 34144 48654 34196
rect 48869 34187 48927 34193
rect 48869 34153 48881 34187
rect 48915 34184 48927 34187
rect 52086 34184 52092 34196
rect 48915 34156 52092 34184
rect 48915 34153 48927 34156
rect 48869 34147 48927 34153
rect 52086 34144 52092 34156
rect 52144 34144 52150 34196
rect 57698 34184 57704 34196
rect 57659 34156 57704 34184
rect 57698 34144 57704 34156
rect 57756 34144 57762 34196
rect 31726 34088 33364 34116
rect 44637 34119 44695 34125
rect 44637 34085 44649 34119
rect 44683 34116 44695 34119
rect 45554 34116 45560 34128
rect 44683 34088 45560 34116
rect 44683 34085 44695 34088
rect 44637 34079 44695 34085
rect 45554 34076 45560 34088
rect 45612 34076 45618 34128
rect 50614 34116 50620 34128
rect 45756 34088 50620 34116
rect 29730 34008 29736 34060
rect 29788 34048 29794 34060
rect 31481 34051 31539 34057
rect 31481 34048 31493 34051
rect 29788 34020 31493 34048
rect 29788 34008 29794 34020
rect 31481 34017 31493 34020
rect 31527 34048 31539 34051
rect 33413 34051 33471 34057
rect 31527 34020 32352 34048
rect 31527 34017 31539 34020
rect 31481 34011 31539 34017
rect 28997 33983 29055 33989
rect 28997 33949 29009 33983
rect 29043 33980 29055 33983
rect 29178 33980 29184 33992
rect 29043 33952 29184 33980
rect 29043 33949 29055 33952
rect 28997 33943 29055 33949
rect 29178 33940 29184 33952
rect 29236 33940 29242 33992
rect 31662 33940 31668 33992
rect 31720 33980 31726 33992
rect 32033 33983 32091 33989
rect 32033 33980 32045 33983
rect 31720 33952 32045 33980
rect 31720 33940 31726 33952
rect 32033 33949 32045 33952
rect 32079 33949 32091 33983
rect 32033 33943 32091 33949
rect 27614 33912 27620 33924
rect 27527 33884 27620 33912
rect 27614 33872 27620 33884
rect 27672 33912 27678 33924
rect 28169 33915 28227 33921
rect 28169 33912 28181 33915
rect 27672 33884 28181 33912
rect 27672 33872 27678 33884
rect 28169 33881 28181 33884
rect 28215 33912 28227 33915
rect 28902 33912 28908 33924
rect 28215 33884 28908 33912
rect 28215 33881 28227 33884
rect 28169 33875 28227 33881
rect 28902 33872 28908 33884
rect 28960 33872 28966 33924
rect 30558 33872 30564 33924
rect 30616 33872 30622 33924
rect 32324 33844 32352 34020
rect 33413 34017 33425 34051
rect 33459 34048 33471 34051
rect 34330 34048 34336 34060
rect 33459 34020 34336 34048
rect 33459 34017 33471 34020
rect 33413 34011 33471 34017
rect 34330 34008 34336 34020
rect 34388 34008 34394 34060
rect 34885 34051 34943 34057
rect 34885 34017 34897 34051
rect 34931 34017 34943 34051
rect 34885 34011 34943 34017
rect 35161 34051 35219 34057
rect 35161 34017 35173 34051
rect 35207 34048 35219 34051
rect 36538 34048 36544 34060
rect 35207 34020 36544 34048
rect 35207 34017 35219 34020
rect 35161 34011 35219 34017
rect 32401 33983 32459 33989
rect 32401 33949 32413 33983
rect 32447 33980 32459 33983
rect 33042 33980 33048 33992
rect 32447 33952 33048 33980
rect 32447 33949 32459 33952
rect 32401 33943 32459 33949
rect 33042 33940 33048 33952
rect 33100 33980 33106 33992
rect 33229 33983 33287 33989
rect 33229 33980 33241 33983
rect 33100 33952 33241 33980
rect 33100 33940 33106 33952
rect 33229 33949 33241 33952
rect 33275 33949 33287 33983
rect 33229 33943 33287 33949
rect 33505 33983 33563 33989
rect 33505 33949 33517 33983
rect 33551 33949 33563 33983
rect 33505 33943 33563 33949
rect 33318 33872 33324 33924
rect 33376 33912 33382 33924
rect 33520 33912 33548 33943
rect 33594 33940 33600 33992
rect 33652 33980 33658 33992
rect 33652 33952 33697 33980
rect 33652 33940 33658 33952
rect 33778 33940 33784 33992
rect 33836 33980 33842 33992
rect 33836 33952 33881 33980
rect 33836 33940 33842 33952
rect 33376 33884 33548 33912
rect 33376 33872 33382 33884
rect 34900 33844 34928 34011
rect 36538 34008 36544 34020
rect 36596 34008 36602 34060
rect 37550 34008 37556 34060
rect 37608 34048 37614 34060
rect 37645 34051 37703 34057
rect 37645 34048 37657 34051
rect 37608 34020 37657 34048
rect 37608 34008 37614 34020
rect 37645 34017 37657 34020
rect 37691 34017 37703 34051
rect 37645 34011 37703 34017
rect 38654 34008 38660 34060
rect 38712 34048 38718 34060
rect 38712 34020 39344 34048
rect 38712 34008 38718 34020
rect 39316 33989 39344 34020
rect 40218 34008 40224 34060
rect 40276 34048 40282 34060
rect 40313 34051 40371 34057
rect 40313 34048 40325 34051
rect 40276 34020 40325 34048
rect 40276 34008 40282 34020
rect 40313 34017 40325 34020
rect 40359 34017 40371 34051
rect 40313 34011 40371 34017
rect 41690 34008 41696 34060
rect 41748 34048 41754 34060
rect 42061 34051 42119 34057
rect 42061 34048 42073 34051
rect 41748 34020 42073 34048
rect 41748 34008 41754 34020
rect 42061 34017 42073 34020
rect 42107 34017 42119 34051
rect 42334 34048 42340 34060
rect 42295 34020 42340 34048
rect 42061 34011 42119 34017
rect 42334 34008 42340 34020
rect 42392 34008 42398 34060
rect 42978 34048 42984 34060
rect 42812 34020 42984 34048
rect 42812 33989 42840 34020
rect 42978 34008 42984 34020
rect 43036 34048 43042 34060
rect 43622 34048 43628 34060
rect 43036 34020 43628 34048
rect 43036 34008 43042 34020
rect 43622 34008 43628 34020
rect 43680 34008 43686 34060
rect 44174 34048 44180 34060
rect 44135 34020 44180 34048
rect 44174 34008 44180 34020
rect 44232 34008 44238 34060
rect 37461 33983 37519 33989
rect 37461 33949 37473 33983
rect 37507 33980 37519 33983
rect 39301 33983 39359 33989
rect 37507 33952 39252 33980
rect 37507 33949 37519 33952
rect 37461 33943 37519 33949
rect 36170 33872 36176 33924
rect 36228 33872 36234 33924
rect 37553 33915 37611 33921
rect 37553 33881 37565 33915
rect 37599 33912 37611 33915
rect 37642 33912 37648 33924
rect 37599 33884 37648 33912
rect 37599 33881 37611 33884
rect 37553 33875 37611 33881
rect 37642 33872 37648 33884
rect 37700 33872 37706 33924
rect 37826 33872 37832 33924
rect 37884 33912 37890 33924
rect 38010 33912 38016 33924
rect 37884 33884 38016 33912
rect 37884 33872 37890 33884
rect 38010 33872 38016 33884
rect 38068 33912 38074 33924
rect 38381 33915 38439 33921
rect 38381 33912 38393 33915
rect 38068 33884 38393 33912
rect 38068 33872 38074 33884
rect 38381 33881 38393 33884
rect 38427 33881 38439 33915
rect 38381 33875 38439 33881
rect 38749 33915 38807 33921
rect 38749 33881 38761 33915
rect 38795 33912 38807 33915
rect 38838 33912 38844 33924
rect 38795 33884 38844 33912
rect 38795 33881 38807 33884
rect 38749 33875 38807 33881
rect 38838 33872 38844 33884
rect 38896 33872 38902 33924
rect 37090 33844 37096 33856
rect 32324 33816 34928 33844
rect 37051 33816 37096 33844
rect 37090 33804 37096 33816
rect 37148 33804 37154 33856
rect 39224 33844 39252 33952
rect 39301 33949 39313 33983
rect 39347 33949 39359 33983
rect 39301 33943 39359 33949
rect 42797 33983 42855 33989
rect 42797 33949 42809 33983
rect 42843 33949 42855 33983
rect 42797 33943 42855 33949
rect 43073 33983 43131 33989
rect 43073 33949 43085 33983
rect 43119 33980 43131 33983
rect 43162 33980 43168 33992
rect 43119 33952 43168 33980
rect 43119 33949 43131 33952
rect 43073 33943 43131 33949
rect 43162 33940 43168 33952
rect 43220 33940 43226 33992
rect 43346 33940 43352 33992
rect 43404 33980 43410 33992
rect 45756 33989 45784 34088
rect 50614 34076 50620 34088
rect 50672 34076 50678 34128
rect 51626 34076 51632 34128
rect 51684 34116 51690 34128
rect 54202 34116 54208 34128
rect 51684 34088 53144 34116
rect 54163 34088 54208 34116
rect 51684 34076 51690 34088
rect 46382 34008 46388 34060
rect 46440 34048 46446 34060
rect 47213 34051 47271 34057
rect 47213 34048 47225 34051
rect 46440 34020 47225 34048
rect 46440 34008 46446 34020
rect 47213 34017 47225 34020
rect 47259 34017 47271 34051
rect 47213 34011 47271 34017
rect 47949 34051 48007 34057
rect 47949 34017 47961 34051
rect 47995 34048 48007 34051
rect 49970 34048 49976 34060
rect 47995 34020 49976 34048
rect 47995 34017 48007 34020
rect 47949 34011 48007 34017
rect 49970 34008 49976 34020
rect 50028 34008 50034 34060
rect 51000 34020 51948 34048
rect 51000 33992 51028 34020
rect 44269 33983 44327 33989
rect 44269 33980 44281 33983
rect 43404 33952 44281 33980
rect 43404 33940 43410 33952
rect 44269 33949 44281 33952
rect 44315 33949 44327 33983
rect 44269 33943 44327 33949
rect 45741 33983 45799 33989
rect 45741 33949 45753 33983
rect 45787 33949 45799 33983
rect 45741 33943 45799 33949
rect 45830 33940 45836 33992
rect 45888 33980 45894 33992
rect 46017 33983 46075 33989
rect 45888 33952 45933 33980
rect 45888 33940 45894 33952
rect 46017 33949 46029 33983
rect 46063 33980 46075 33983
rect 47121 33983 47179 33989
rect 46063 33952 46704 33980
rect 46063 33949 46075 33952
rect 46017 33943 46075 33949
rect 41966 33912 41972 33924
rect 41630 33884 41972 33912
rect 41966 33872 41972 33884
rect 42024 33872 42030 33924
rect 42058 33872 42064 33924
rect 42116 33912 42122 33924
rect 42610 33912 42616 33924
rect 42116 33884 42616 33912
rect 42116 33872 42122 33884
rect 42610 33872 42616 33884
rect 42668 33912 42674 33924
rect 45189 33915 45247 33921
rect 45189 33912 45201 33915
rect 42668 33884 45201 33912
rect 42668 33872 42674 33884
rect 45189 33881 45201 33884
rect 45235 33881 45247 33915
rect 45189 33875 45247 33881
rect 42794 33844 42800 33856
rect 39224 33816 42800 33844
rect 42794 33804 42800 33816
rect 42852 33804 42858 33856
rect 42889 33847 42947 33853
rect 42889 33813 42901 33847
rect 42935 33844 42947 33847
rect 43254 33844 43260 33856
rect 42935 33816 43260 33844
rect 42935 33813 42947 33816
rect 42889 33807 42947 33813
rect 43254 33804 43260 33816
rect 43312 33804 43318 33856
rect 46198 33844 46204 33856
rect 46159 33816 46204 33844
rect 46198 33804 46204 33816
rect 46256 33804 46262 33856
rect 46676 33853 46704 33952
rect 47121 33949 47133 33983
rect 47167 33980 47179 33983
rect 48682 33980 48688 33992
rect 47167 33952 48688 33980
rect 47167 33949 47179 33952
rect 47121 33943 47179 33949
rect 48682 33940 48688 33952
rect 48740 33940 48746 33992
rect 48774 33940 48780 33992
rect 48832 33980 48838 33992
rect 49421 33983 49479 33989
rect 49421 33980 49433 33983
rect 48832 33952 49433 33980
rect 48832 33940 48838 33952
rect 49421 33949 49433 33952
rect 49467 33949 49479 33983
rect 49602 33980 49608 33992
rect 49563 33952 49608 33980
rect 49421 33943 49479 33949
rect 49602 33940 49608 33952
rect 49660 33940 49666 33992
rect 50982 33980 50988 33992
rect 50943 33952 50988 33980
rect 50982 33940 50988 33952
rect 51040 33940 51046 33992
rect 51920 33989 51948 34020
rect 51077 33983 51135 33989
rect 51077 33949 51089 33983
rect 51123 33949 51135 33983
rect 51077 33943 51135 33949
rect 51905 33983 51963 33989
rect 51905 33949 51917 33983
rect 51951 33949 51963 33983
rect 52086 33980 52092 33992
rect 52047 33952 52092 33980
rect 51905 33943 51963 33949
rect 47029 33915 47087 33921
rect 47029 33881 47041 33915
rect 47075 33912 47087 33915
rect 47762 33912 47768 33924
rect 47075 33884 47768 33912
rect 47075 33881 47087 33884
rect 47029 33875 47087 33881
rect 47762 33872 47768 33884
rect 47820 33872 47826 33924
rect 48409 33915 48467 33921
rect 48409 33881 48421 33915
rect 48455 33912 48467 33915
rect 48590 33912 48596 33924
rect 48455 33884 48596 33912
rect 48455 33881 48467 33884
rect 48409 33875 48467 33881
rect 48590 33872 48596 33884
rect 48648 33912 48654 33924
rect 49326 33912 49332 33924
rect 48648 33884 49332 33912
rect 48648 33872 48654 33884
rect 49326 33872 49332 33884
rect 49384 33912 49390 33924
rect 49513 33915 49571 33921
rect 49513 33912 49525 33915
rect 49384 33884 49525 33912
rect 49384 33872 49390 33884
rect 49513 33881 49525 33884
rect 49559 33881 49571 33915
rect 49513 33875 49571 33881
rect 49694 33872 49700 33924
rect 49752 33912 49758 33924
rect 51092 33912 51120 33943
rect 52086 33940 52092 33952
rect 52144 33940 52150 33992
rect 51350 33912 51356 33924
rect 49752 33884 50936 33912
rect 51092 33884 51356 33912
rect 49752 33872 49758 33884
rect 46661 33847 46719 33853
rect 46661 33813 46673 33847
rect 46707 33813 46719 33847
rect 46661 33807 46719 33813
rect 48314 33804 48320 33856
rect 48372 33844 48378 33856
rect 48501 33847 48559 33853
rect 48501 33844 48513 33847
rect 48372 33816 48513 33844
rect 48372 33804 48378 33816
rect 48501 33813 48513 33816
rect 48547 33813 48559 33847
rect 48501 33807 48559 33813
rect 50246 33804 50252 33856
rect 50304 33844 50310 33856
rect 50801 33847 50859 33853
rect 50801 33844 50813 33847
rect 50304 33816 50813 33844
rect 50304 33804 50310 33816
rect 50801 33813 50813 33816
rect 50847 33813 50859 33847
rect 50908 33844 50936 33884
rect 51350 33872 51356 33884
rect 51408 33912 51414 33924
rect 52104 33912 52132 33940
rect 51408 33884 52132 33912
rect 51408 33872 51414 33884
rect 51445 33847 51503 33853
rect 51445 33844 51457 33847
rect 50908 33816 51457 33844
rect 50801 33807 50859 33813
rect 51445 33813 51457 33816
rect 51491 33844 51503 33847
rect 51626 33844 51632 33856
rect 51491 33816 51632 33844
rect 51491 33813 51503 33816
rect 51445 33807 51503 33813
rect 51626 33804 51632 33816
rect 51684 33804 51690 33856
rect 51994 33844 52000 33856
rect 51955 33816 52000 33844
rect 51994 33804 52000 33816
rect 52052 33804 52058 33856
rect 53006 33844 53012 33856
rect 52967 33816 53012 33844
rect 53006 33804 53012 33816
rect 53064 33804 53070 33856
rect 53116 33844 53144 34088
rect 54202 34076 54208 34088
rect 54260 34076 54266 34128
rect 55769 34051 55827 34057
rect 55769 34048 55781 34051
rect 53208 34020 55781 34048
rect 53208 33989 53236 34020
rect 55769 34017 55781 34020
rect 55815 34017 55827 34051
rect 55769 34011 55827 34017
rect 53193 33983 53251 33989
rect 53193 33949 53205 33983
rect 53239 33949 53251 33983
rect 53193 33943 53251 33949
rect 53377 33983 53435 33989
rect 53377 33949 53389 33983
rect 53423 33949 53435 33983
rect 53377 33943 53435 33949
rect 53469 33983 53527 33989
rect 53469 33949 53481 33983
rect 53515 33980 53527 33983
rect 54018 33980 54024 33992
rect 53515 33952 54024 33980
rect 53515 33949 53527 33952
rect 53469 33943 53527 33949
rect 53392 33912 53420 33943
rect 54018 33940 54024 33952
rect 54076 33940 54082 33992
rect 54478 33980 54484 33992
rect 54439 33952 54484 33980
rect 54478 33940 54484 33952
rect 54536 33940 54542 33992
rect 55950 33980 55956 33992
rect 55911 33952 55956 33980
rect 55950 33940 55956 33952
rect 56008 33940 56014 33992
rect 56042 33940 56048 33992
rect 56100 33980 56106 33992
rect 56226 33980 56232 33992
rect 56100 33952 56145 33980
rect 56187 33952 56232 33980
rect 56100 33940 56106 33952
rect 56226 33940 56232 33952
rect 56284 33940 56290 33992
rect 56321 33983 56379 33989
rect 56321 33949 56333 33983
rect 56367 33980 56379 33983
rect 56962 33980 56968 33992
rect 56367 33952 56968 33980
rect 56367 33949 56379 33952
rect 56321 33943 56379 33949
rect 56962 33940 56968 33952
rect 57020 33940 57026 33992
rect 53558 33912 53564 33924
rect 53392 33884 53564 33912
rect 53558 33872 53564 33884
rect 53616 33872 53622 33924
rect 54205 33915 54263 33921
rect 54205 33881 54217 33915
rect 54251 33912 54263 33915
rect 55766 33912 55772 33924
rect 54251 33884 55772 33912
rect 54251 33881 54263 33884
rect 54205 33875 54263 33881
rect 54220 33844 54248 33875
rect 55766 33872 55772 33884
rect 55824 33872 55830 33924
rect 55858 33872 55864 33924
rect 55916 33912 55922 33924
rect 56244 33912 56272 33940
rect 55916 33884 56272 33912
rect 55916 33872 55922 33884
rect 56594 33872 56600 33924
rect 56652 33912 56658 33924
rect 57609 33915 57667 33921
rect 57609 33912 57621 33915
rect 56652 33884 57621 33912
rect 56652 33872 56658 33884
rect 57609 33881 57621 33884
rect 57655 33881 57667 33915
rect 57609 33875 57667 33881
rect 54386 33844 54392 33856
rect 53116 33816 54248 33844
rect 54347 33816 54392 33844
rect 54386 33804 54392 33816
rect 54444 33804 54450 33856
rect 56778 33844 56784 33856
rect 56739 33816 56784 33844
rect 56778 33804 56784 33816
rect 56836 33804 56842 33856
rect 1104 33754 58880 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 58880 33754
rect 1104 33680 58880 33702
rect 31481 33643 31539 33649
rect 31481 33609 31493 33643
rect 31527 33609 31539 33643
rect 31481 33603 31539 33609
rect 33413 33643 33471 33649
rect 33413 33609 33425 33643
rect 33459 33640 33471 33643
rect 33594 33640 33600 33652
rect 33459 33612 33600 33640
rect 33459 33609 33471 33612
rect 33413 33603 33471 33609
rect 31018 33532 31024 33584
rect 31076 33532 31082 33584
rect 31496 33572 31524 33603
rect 33594 33600 33600 33612
rect 33652 33600 33658 33652
rect 34698 33600 34704 33652
rect 34756 33640 34762 33652
rect 35345 33643 35403 33649
rect 35345 33640 35357 33643
rect 34756 33612 35357 33640
rect 34756 33600 34762 33612
rect 35345 33609 35357 33612
rect 35391 33609 35403 33643
rect 35345 33603 35403 33609
rect 38838 33600 38844 33652
rect 38896 33640 38902 33652
rect 41966 33640 41972 33652
rect 38896 33612 39988 33640
rect 41927 33612 41972 33640
rect 38896 33600 38902 33612
rect 31754 33572 31760 33584
rect 31496 33544 31760 33572
rect 31754 33532 31760 33544
rect 31812 33572 31818 33584
rect 32401 33575 32459 33581
rect 32401 33572 32413 33575
rect 31812 33544 32413 33572
rect 31812 33532 31818 33544
rect 32401 33541 32413 33544
rect 32447 33541 32459 33575
rect 32401 33535 32459 33541
rect 32769 33575 32827 33581
rect 32769 33541 32781 33575
rect 32815 33572 32827 33575
rect 33778 33572 33784 33584
rect 32815 33544 33784 33572
rect 32815 33541 32827 33544
rect 32769 33535 32827 33541
rect 33778 33532 33784 33544
rect 33836 33572 33842 33584
rect 33836 33544 36584 33572
rect 33836 33532 33842 33544
rect 28074 33464 28080 33516
rect 28132 33504 28138 33516
rect 29730 33504 29736 33516
rect 28132 33476 29736 33504
rect 28132 33464 28138 33476
rect 29730 33464 29736 33476
rect 29788 33464 29794 33516
rect 33226 33504 33232 33516
rect 33187 33476 33232 33504
rect 33226 33464 33232 33476
rect 33284 33464 33290 33516
rect 33413 33507 33471 33513
rect 33413 33473 33425 33507
rect 33459 33473 33471 33507
rect 34698 33504 34704 33516
rect 34659 33476 34704 33504
rect 33413 33467 33471 33473
rect 30009 33439 30067 33445
rect 30009 33405 30021 33439
rect 30055 33436 30067 33439
rect 30055 33408 31754 33436
rect 30055 33405 30067 33408
rect 30009 33399 30067 33405
rect 28721 33303 28779 33309
rect 28721 33269 28733 33303
rect 28767 33300 28779 33303
rect 29178 33300 29184 33312
rect 28767 33272 29184 33300
rect 28767 33269 28779 33272
rect 28721 33263 28779 33269
rect 29178 33260 29184 33272
rect 29236 33260 29242 33312
rect 31726 33300 31754 33408
rect 33042 33396 33048 33448
rect 33100 33436 33106 33448
rect 33428 33436 33456 33467
rect 34698 33464 34704 33476
rect 34756 33504 34762 33516
rect 36556 33513 36584 33544
rect 38930 33532 38936 33584
rect 38988 33532 38994 33584
rect 39960 33581 39988 33612
rect 41966 33600 41972 33612
rect 42024 33600 42030 33652
rect 47210 33600 47216 33652
rect 47268 33640 47274 33652
rect 49694 33640 49700 33652
rect 47268 33612 49700 33640
rect 47268 33600 47274 33612
rect 49694 33600 49700 33612
rect 49752 33600 49758 33652
rect 53558 33640 53564 33652
rect 50908 33612 53052 33640
rect 53519 33612 53564 33640
rect 39945 33575 40003 33581
rect 39945 33541 39957 33575
rect 39991 33572 40003 33575
rect 39991 33544 43668 33572
rect 39991 33541 40003 33544
rect 39945 33535 40003 33541
rect 35161 33507 35219 33513
rect 35161 33504 35173 33507
rect 34756 33476 35173 33504
rect 34756 33464 34762 33476
rect 35161 33473 35173 33476
rect 35207 33473 35219 33507
rect 35161 33467 35219 33473
rect 36541 33507 36599 33513
rect 36541 33473 36553 33507
rect 36587 33504 36599 33507
rect 37274 33504 37280 33516
rect 36587 33476 37280 33504
rect 36587 33473 36599 33476
rect 36541 33467 36599 33473
rect 37274 33464 37280 33476
rect 37332 33504 37338 33516
rect 37734 33504 37740 33516
rect 37332 33476 37740 33504
rect 37332 33464 37338 33476
rect 37734 33464 37740 33476
rect 37792 33464 37798 33516
rect 39482 33464 39488 33516
rect 39540 33504 39546 33516
rect 41417 33507 41475 33513
rect 41417 33504 41429 33507
rect 39540 33476 41429 33504
rect 39540 33464 39546 33476
rect 41417 33473 41429 33476
rect 41463 33473 41475 33507
rect 42058 33504 42064 33516
rect 42019 33476 42064 33504
rect 41417 33467 41475 33473
rect 42058 33464 42064 33476
rect 42116 33464 42122 33516
rect 42981 33507 43039 33513
rect 42981 33473 42993 33507
rect 43027 33504 43039 33507
rect 43346 33504 43352 33516
rect 43027 33476 43352 33504
rect 43027 33473 43039 33476
rect 42981 33467 43039 33473
rect 43346 33464 43352 33476
rect 43404 33504 43410 33516
rect 43640 33513 43668 33544
rect 45462 33532 45468 33584
rect 45520 33572 45526 33584
rect 50908 33572 50936 33612
rect 51994 33572 52000 33584
rect 45520 33544 50936 33572
rect 51046 33544 52000 33572
rect 45520 33532 45526 33544
rect 43533 33507 43591 33513
rect 43533 33504 43545 33507
rect 43404 33476 43545 33504
rect 43404 33464 43410 33476
rect 43533 33473 43545 33476
rect 43579 33473 43591 33507
rect 43533 33467 43591 33473
rect 43625 33507 43683 33513
rect 43625 33473 43637 33507
rect 43671 33504 43683 33507
rect 43898 33504 43904 33516
rect 43671 33476 43904 33504
rect 43671 33473 43683 33476
rect 43625 33467 43683 33473
rect 43898 33464 43904 33476
rect 43956 33464 43962 33516
rect 44542 33504 44548 33516
rect 44503 33476 44548 33504
rect 44542 33464 44548 33476
rect 44600 33464 44606 33516
rect 44634 33464 44640 33516
rect 44692 33504 44698 33516
rect 44821 33507 44879 33513
rect 44692 33476 44737 33504
rect 44692 33464 44698 33476
rect 44821 33473 44833 33507
rect 44867 33473 44879 33507
rect 46014 33504 46020 33516
rect 45975 33476 46020 33504
rect 44821 33467 44879 33473
rect 33100 33408 33456 33436
rect 36633 33439 36691 33445
rect 33100 33396 33106 33408
rect 36633 33405 36645 33439
rect 36679 33436 36691 33439
rect 37090 33436 37096 33448
rect 36679 33408 37096 33436
rect 36679 33405 36691 33408
rect 36633 33399 36691 33405
rect 37090 33396 37096 33408
rect 37148 33396 37154 33448
rect 37921 33439 37979 33445
rect 37921 33405 37933 33439
rect 37967 33405 37979 33439
rect 38194 33436 38200 33448
rect 38155 33408 38200 33436
rect 37921 33399 37979 33405
rect 34440 33340 35388 33368
rect 34440 33300 34468 33340
rect 31726 33272 34468 33300
rect 34517 33303 34575 33309
rect 34517 33269 34529 33303
rect 34563 33300 34575 33303
rect 34606 33300 34612 33312
rect 34563 33272 34612 33300
rect 34563 33269 34575 33272
rect 34517 33263 34575 33269
rect 34606 33260 34612 33272
rect 34664 33260 34670 33312
rect 35360 33300 35388 33340
rect 35434 33328 35440 33380
rect 35492 33368 35498 33380
rect 37936 33368 37964 33399
rect 38194 33396 38200 33408
rect 38252 33396 38258 33448
rect 42702 33436 42708 33448
rect 42663 33408 42708 33436
rect 42702 33396 42708 33408
rect 42760 33396 42766 33448
rect 43162 33396 43168 33448
rect 43220 33436 43226 33448
rect 44836 33436 44864 33467
rect 46014 33464 46020 33476
rect 46072 33464 46078 33516
rect 48222 33504 48228 33516
rect 48183 33476 48228 33504
rect 48222 33464 48228 33476
rect 48280 33464 48286 33516
rect 48498 33504 48504 33516
rect 48459 33476 48504 33504
rect 48498 33464 48504 33476
rect 48556 33464 48562 33516
rect 48682 33504 48688 33516
rect 48643 33476 48688 33504
rect 48682 33464 48688 33476
rect 48740 33464 48746 33516
rect 49970 33504 49976 33516
rect 49931 33476 49976 33504
rect 49970 33464 49976 33476
rect 50028 33464 50034 33516
rect 50246 33504 50252 33516
rect 50207 33476 50252 33504
rect 50246 33464 50252 33476
rect 50304 33464 50310 33516
rect 50433 33507 50491 33513
rect 50433 33473 50445 33507
rect 50479 33504 50491 33507
rect 51046 33504 51074 33544
rect 51994 33532 52000 33544
rect 52052 33532 52058 33584
rect 52454 33572 52460 33584
rect 52196 33544 52460 33572
rect 51350 33504 51356 33516
rect 50479 33476 51074 33504
rect 51311 33476 51356 33504
rect 50479 33473 50491 33476
rect 50433 33467 50491 33473
rect 51350 33464 51356 33476
rect 51408 33464 51414 33516
rect 52196 33513 52224 33544
rect 52454 33532 52460 33544
rect 52512 33532 52518 33584
rect 53024 33572 53052 33612
rect 53558 33600 53564 33612
rect 53616 33600 53622 33652
rect 54018 33640 54024 33652
rect 53979 33612 54024 33640
rect 54018 33600 54024 33612
rect 54076 33600 54082 33652
rect 57054 33600 57060 33652
rect 57112 33640 57118 33652
rect 57422 33640 57428 33652
rect 57112 33612 57428 33640
rect 57112 33600 57118 33612
rect 57422 33600 57428 33612
rect 57480 33600 57486 33652
rect 53650 33572 53656 33584
rect 53024 33544 53656 33572
rect 53650 33532 53656 33544
rect 53708 33532 53714 33584
rect 54478 33572 54484 33584
rect 54404 33544 54484 33572
rect 52181 33507 52239 33513
rect 52181 33473 52193 33507
rect 52227 33473 52239 33507
rect 52362 33504 52368 33516
rect 52323 33476 52368 33504
rect 52181 33467 52239 33473
rect 52362 33464 52368 33476
rect 52420 33464 52426 33516
rect 53190 33504 53196 33516
rect 52932 33476 53196 33504
rect 48406 33436 48412 33448
rect 43220 33408 44864 33436
rect 48367 33408 48412 33436
rect 43220 33396 43226 33408
rect 48406 33396 48412 33408
rect 48464 33396 48470 33448
rect 49786 33396 49792 33448
rect 49844 33436 49850 33448
rect 50157 33439 50215 33445
rect 50157 33436 50169 33439
rect 49844 33408 50169 33436
rect 49844 33396 49850 33408
rect 50157 33405 50169 33408
rect 50203 33405 50215 33439
rect 50982 33436 50988 33448
rect 50943 33408 50988 33436
rect 50157 33399 50215 33405
rect 50982 33396 50988 33408
rect 51040 33396 51046 33448
rect 51074 33396 51080 33448
rect 51132 33436 51138 33448
rect 51261 33439 51319 33445
rect 51261 33436 51273 33439
rect 51132 33408 51273 33436
rect 51132 33396 51138 33408
rect 51261 33405 51273 33408
rect 51307 33405 51319 33439
rect 52932 33436 52960 33476
rect 53190 33464 53196 33476
rect 53248 33464 53254 33516
rect 53374 33504 53380 33516
rect 53335 33476 53380 33504
rect 53374 33464 53380 33476
rect 53432 33464 53438 33516
rect 54202 33504 54208 33516
rect 54163 33476 54208 33504
rect 54202 33464 54208 33476
rect 54260 33464 54266 33516
rect 54404 33513 54432 33544
rect 54478 33532 54484 33544
rect 54536 33532 54542 33584
rect 54389 33507 54447 33513
rect 54389 33473 54401 33507
rect 54435 33473 54447 33507
rect 54389 33467 54447 33473
rect 56594 33464 56600 33516
rect 56652 33504 56658 33516
rect 57057 33507 57115 33513
rect 57057 33504 57069 33507
rect 56652 33476 57069 33504
rect 56652 33464 56658 33476
rect 57057 33473 57069 33476
rect 57103 33473 57115 33507
rect 57057 33467 57115 33473
rect 57514 33464 57520 33516
rect 57572 33504 57578 33516
rect 57572 33476 57617 33504
rect 57572 33464 57578 33476
rect 53098 33436 53104 33448
rect 51261 33399 51319 33405
rect 52197 33408 52960 33436
rect 53059 33408 53104 33436
rect 35492 33340 37964 33368
rect 35492 33328 35498 33340
rect 36722 33300 36728 33312
rect 35360 33272 36728 33300
rect 36722 33260 36728 33272
rect 36780 33260 36786 33312
rect 36817 33303 36875 33309
rect 36817 33269 36829 33303
rect 36863 33300 36875 33303
rect 37090 33300 37096 33312
rect 36863 33272 37096 33300
rect 36863 33269 36875 33272
rect 36817 33263 36875 33269
rect 37090 33260 37096 33272
rect 37148 33260 37154 33312
rect 37936 33300 37964 33340
rect 42797 33371 42855 33377
rect 42797 33337 42809 33371
rect 42843 33368 42855 33371
rect 42978 33368 42984 33380
rect 42843 33340 42984 33368
rect 42843 33337 42855 33340
rect 42797 33331 42855 33337
rect 42978 33328 42984 33340
rect 43036 33328 43042 33380
rect 45005 33371 45063 33377
rect 45005 33337 45017 33371
rect 45051 33368 45063 33371
rect 46382 33368 46388 33380
rect 45051 33340 46388 33368
rect 45051 33337 45063 33340
rect 45005 33331 45063 33337
rect 46382 33328 46388 33340
rect 46440 33328 46446 33380
rect 47854 33328 47860 33380
rect 47912 33368 47918 33380
rect 48593 33371 48651 33377
rect 48593 33368 48605 33371
rect 47912 33340 48605 33368
rect 47912 33328 47918 33340
rect 48593 33337 48605 33340
rect 48639 33337 48651 33371
rect 50062 33368 50068 33380
rect 50023 33340 50068 33368
rect 48593 33331 48651 33337
rect 50062 33328 50068 33340
rect 50120 33328 50126 33380
rect 52197 33368 52225 33408
rect 53098 33396 53104 33408
rect 53156 33396 53162 33448
rect 53285 33439 53343 33445
rect 53285 33405 53297 33439
rect 53331 33405 53343 33439
rect 54478 33436 54484 33448
rect 54439 33408 54484 33436
rect 53285 33399 53343 33405
rect 51046 33340 52225 33368
rect 52273 33371 52331 33377
rect 38286 33300 38292 33312
rect 37936 33272 38292 33300
rect 38286 33260 38292 33272
rect 38344 33300 38350 33312
rect 40405 33303 40463 33309
rect 40405 33300 40417 33303
rect 38344 33272 40417 33300
rect 38344 33260 38350 33272
rect 40405 33269 40417 33272
rect 40451 33269 40463 33303
rect 40405 33263 40463 33269
rect 41325 33303 41383 33309
rect 41325 33269 41337 33303
rect 41371 33300 41383 33303
rect 41414 33300 41420 33312
rect 41371 33272 41420 33300
rect 41371 33269 41383 33272
rect 41325 33263 41383 33269
rect 41414 33260 41420 33272
rect 41472 33260 41478 33312
rect 41506 33260 41512 33312
rect 41564 33300 41570 33312
rect 42889 33303 42947 33309
rect 42889 33300 42901 33303
rect 41564 33272 42901 33300
rect 41564 33260 41570 33272
rect 42889 33269 42901 33272
rect 42935 33300 42947 33303
rect 45186 33300 45192 33312
rect 42935 33272 45192 33300
rect 42935 33269 42947 33272
rect 42889 33263 42947 33269
rect 45186 33260 45192 33272
rect 45244 33260 45250 33312
rect 45922 33260 45928 33312
rect 45980 33300 45986 33312
rect 46109 33303 46167 33309
rect 46109 33300 46121 33303
rect 45980 33272 46121 33300
rect 45980 33260 45986 33272
rect 46109 33269 46121 33272
rect 46155 33269 46167 33303
rect 46109 33263 46167 33269
rect 46937 33303 46995 33309
rect 46937 33269 46949 33303
rect 46983 33300 46995 33303
rect 47026 33300 47032 33312
rect 46983 33272 47032 33300
rect 46983 33269 46995 33272
rect 46937 33263 46995 33269
rect 47026 33260 47032 33272
rect 47084 33260 47090 33312
rect 48869 33303 48927 33309
rect 48869 33269 48881 33303
rect 48915 33300 48927 33303
rect 49602 33300 49608 33312
rect 48915 33272 49608 33300
rect 48915 33269 48927 33272
rect 48869 33263 48927 33269
rect 49602 33260 49608 33272
rect 49660 33260 49666 33312
rect 49694 33260 49700 33312
rect 49752 33300 49758 33312
rect 49789 33303 49847 33309
rect 49789 33300 49801 33303
rect 49752 33272 49801 33300
rect 49752 33260 49758 33272
rect 49789 33269 49801 33272
rect 49835 33269 49847 33303
rect 49789 33263 49847 33269
rect 49970 33260 49976 33312
rect 50028 33300 50034 33312
rect 51046 33300 51074 33340
rect 52273 33337 52285 33371
rect 52319 33368 52331 33371
rect 53300 33368 53328 33399
rect 54478 33396 54484 33408
rect 54536 33396 54542 33448
rect 54938 33396 54944 33448
rect 54996 33436 55002 33448
rect 55493 33439 55551 33445
rect 55493 33436 55505 33439
rect 54996 33408 55505 33436
rect 54996 33396 55002 33408
rect 55493 33405 55505 33408
rect 55539 33436 55551 33439
rect 56778 33436 56784 33448
rect 55539 33408 56784 33436
rect 55539 33405 55551 33408
rect 55493 33399 55551 33405
rect 56778 33396 56784 33408
rect 56836 33396 56842 33448
rect 57882 33396 57888 33448
rect 57940 33396 57946 33448
rect 57974 33396 57980 33448
rect 58032 33436 58038 33448
rect 58069 33439 58127 33445
rect 58069 33436 58081 33439
rect 58032 33408 58081 33436
rect 58032 33396 58038 33408
rect 58069 33405 58081 33408
rect 58115 33405 58127 33439
rect 58069 33399 58127 33405
rect 52319 33340 53328 33368
rect 52319 33337 52331 33340
rect 52273 33331 52331 33337
rect 54110 33328 54116 33380
rect 54168 33368 54174 33380
rect 55398 33368 55404 33380
rect 54168 33340 55404 33368
rect 54168 33328 54174 33340
rect 55398 33328 55404 33340
rect 55456 33368 55462 33380
rect 56045 33371 56103 33377
rect 56045 33368 56057 33371
rect 55456 33340 56057 33368
rect 55456 33328 55462 33340
rect 56045 33337 56057 33340
rect 56091 33337 56103 33371
rect 56045 33331 56103 33337
rect 56686 33328 56692 33380
rect 56744 33368 56750 33380
rect 57900 33368 57928 33396
rect 56744 33340 57928 33368
rect 56744 33328 56750 33340
rect 50028 33272 51074 33300
rect 50028 33260 50034 33272
rect 53650 33260 53656 33312
rect 53708 33300 53714 33312
rect 54941 33303 54999 33309
rect 54941 33300 54953 33303
rect 53708 33272 54953 33300
rect 53708 33260 53714 33272
rect 54941 33269 54953 33272
rect 54987 33269 54999 33303
rect 54941 33263 54999 33269
rect 57241 33303 57299 33309
rect 57241 33269 57253 33303
rect 57287 33300 57299 33303
rect 57974 33300 57980 33312
rect 57287 33272 57980 33300
rect 57287 33269 57299 33272
rect 57241 33263 57299 33269
rect 57974 33260 57980 33272
rect 58032 33260 58038 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 29178 33096 29184 33108
rect 29139 33068 29184 33096
rect 29178 33056 29184 33068
rect 29236 33056 29242 33108
rect 30558 33096 30564 33108
rect 30519 33068 30564 33096
rect 30558 33056 30564 33068
rect 30616 33056 30622 33108
rect 33045 33099 33103 33105
rect 33045 33065 33057 33099
rect 33091 33096 33103 33099
rect 34146 33096 34152 33108
rect 33091 33068 34152 33096
rect 33091 33065 33103 33068
rect 33045 33059 33103 33065
rect 34146 33056 34152 33068
rect 34204 33056 34210 33108
rect 34606 33056 34612 33108
rect 34664 33096 34670 33108
rect 35342 33096 35348 33108
rect 34664 33068 35348 33096
rect 34664 33056 34670 33068
rect 35342 33056 35348 33068
rect 35400 33096 35406 33108
rect 36538 33096 36544 33108
rect 35400 33068 36216 33096
rect 36499 33068 36544 33096
rect 35400 33056 35406 33068
rect 36081 33031 36139 33037
rect 36081 32997 36093 33031
rect 36127 32997 36139 33031
rect 36081 32991 36139 32997
rect 29730 32920 29736 32972
rect 29788 32960 29794 32972
rect 31297 32963 31355 32969
rect 31297 32960 31309 32963
rect 29788 32932 31309 32960
rect 29788 32920 29794 32932
rect 31297 32929 31309 32932
rect 31343 32929 31355 32963
rect 31297 32923 31355 32929
rect 35437 32963 35495 32969
rect 35437 32929 35449 32963
rect 35483 32929 35495 32963
rect 35437 32923 35495 32929
rect 29178 32852 29184 32904
rect 29236 32892 29242 32904
rect 29917 32895 29975 32901
rect 29917 32892 29929 32895
rect 29236 32864 29929 32892
rect 29236 32852 29242 32864
rect 29917 32861 29929 32864
rect 29963 32892 29975 32895
rect 30282 32892 30288 32904
rect 29963 32864 30288 32892
rect 29963 32861 29975 32864
rect 29917 32855 29975 32861
rect 30282 32852 30288 32864
rect 30340 32892 30346 32904
rect 30653 32895 30711 32901
rect 30653 32892 30665 32895
rect 30340 32864 30665 32892
rect 30340 32852 30346 32864
rect 30653 32861 30665 32864
rect 30699 32861 30711 32895
rect 30653 32855 30711 32861
rect 32858 32852 32864 32904
rect 32916 32892 32922 32904
rect 33781 32895 33839 32901
rect 33781 32892 33793 32895
rect 32916 32864 33793 32892
rect 32916 32852 32922 32864
rect 33781 32861 33793 32864
rect 33827 32861 33839 32895
rect 33781 32855 33839 32861
rect 34790 32852 34796 32904
rect 34848 32892 34854 32904
rect 35452 32892 35480 32923
rect 34848 32864 35480 32892
rect 35713 32895 35771 32901
rect 34848 32852 34854 32864
rect 35713 32861 35725 32895
rect 35759 32892 35771 32895
rect 36096 32892 36124 32991
rect 36188 32960 36216 33068
rect 36538 33056 36544 33068
rect 36596 33056 36602 33108
rect 38930 33056 38936 33108
rect 38988 33096 38994 33108
rect 39025 33099 39083 33105
rect 39025 33096 39037 33099
rect 38988 33068 39037 33096
rect 38988 33056 38994 33068
rect 39025 33065 39037 33068
rect 39071 33065 39083 33099
rect 41874 33096 41880 33108
rect 39025 33059 39083 33065
rect 40236 33068 41736 33096
rect 41835 33068 41880 33096
rect 36722 32988 36728 33040
rect 36780 33028 36786 33040
rect 37185 33031 37243 33037
rect 37185 33028 37197 33031
rect 36780 33000 37197 33028
rect 36780 32988 36786 33000
rect 37185 32997 37197 33000
rect 37231 32997 37243 33031
rect 40236 33028 40264 33068
rect 37185 32991 37243 32997
rect 37292 33000 40264 33028
rect 36906 32960 36912 32972
rect 36188 32932 36912 32960
rect 36906 32920 36912 32932
rect 36964 32920 36970 32972
rect 37292 32960 37320 33000
rect 39850 32960 39856 32972
rect 37200 32932 37320 32960
rect 37476 32932 39856 32960
rect 37200 32904 37228 32932
rect 36725 32895 36783 32901
rect 36725 32892 36737 32895
rect 35759 32864 36032 32892
rect 36096 32864 36737 32892
rect 35759 32861 35771 32864
rect 35713 32855 35771 32861
rect 31570 32824 31576 32836
rect 31531 32796 31576 32824
rect 31570 32784 31576 32796
rect 31628 32784 31634 32836
rect 33689 32827 33747 32833
rect 33689 32824 33701 32827
rect 32798 32796 33701 32824
rect 33689 32793 33701 32796
rect 33735 32793 33747 32827
rect 33689 32787 33747 32793
rect 35621 32827 35679 32833
rect 35621 32793 35633 32827
rect 35667 32824 35679 32827
rect 36004 32824 36032 32864
rect 36725 32861 36737 32864
rect 36771 32861 36783 32895
rect 36725 32855 36783 32861
rect 37182 32852 37188 32904
rect 37240 32852 37246 32904
rect 37366 32892 37372 32904
rect 37327 32864 37372 32892
rect 37366 32852 37372 32864
rect 37424 32852 37430 32904
rect 37476 32901 37504 32932
rect 39850 32920 39856 32932
rect 39908 32920 39914 32972
rect 40129 32963 40187 32969
rect 40129 32929 40141 32963
rect 40175 32960 40187 32963
rect 41046 32960 41052 32972
rect 40175 32932 41052 32960
rect 40175 32929 40187 32932
rect 40129 32923 40187 32929
rect 41046 32920 41052 32932
rect 41104 32920 41110 32972
rect 41708 32960 41736 33068
rect 41874 33056 41880 33068
rect 41932 33056 41938 33108
rect 48406 33056 48412 33108
rect 48464 33096 48470 33108
rect 48501 33099 48559 33105
rect 48501 33096 48513 33099
rect 48464 33068 48513 33096
rect 48464 33056 48470 33068
rect 48501 33065 48513 33068
rect 48547 33065 48559 33099
rect 49786 33096 49792 33108
rect 49747 33068 49792 33096
rect 48501 33059 48559 33065
rect 49786 33056 49792 33068
rect 49844 33056 49850 33108
rect 50062 33056 50068 33108
rect 50120 33096 50126 33108
rect 50341 33099 50399 33105
rect 50341 33096 50353 33099
rect 50120 33068 50353 33096
rect 50120 33056 50126 33068
rect 50341 33065 50353 33068
rect 50387 33065 50399 33099
rect 50341 33059 50399 33065
rect 50798 33056 50804 33108
rect 50856 33096 50862 33108
rect 52273 33099 52331 33105
rect 50856 33068 51304 33096
rect 50856 33056 50862 33068
rect 46661 33031 46719 33037
rect 46661 32997 46673 33031
rect 46707 33028 46719 33031
rect 46707 33000 47348 33028
rect 46707 32997 46719 33000
rect 46661 32991 46719 32997
rect 41708 32932 43024 32960
rect 37461 32895 37519 32901
rect 37461 32861 37473 32895
rect 37507 32861 37519 32895
rect 37734 32892 37740 32904
rect 37695 32864 37740 32892
rect 37461 32855 37519 32861
rect 37734 32852 37740 32864
rect 37792 32852 37798 32904
rect 37918 32852 37924 32904
rect 37976 32892 37982 32904
rect 38562 32892 38568 32904
rect 37976 32864 38568 32892
rect 37976 32852 37982 32864
rect 38562 32852 38568 32864
rect 38620 32852 38626 32904
rect 38654 32852 38660 32904
rect 38712 32892 38718 32904
rect 38933 32895 38991 32901
rect 38933 32892 38945 32895
rect 38712 32864 38945 32892
rect 38712 32852 38718 32864
rect 38933 32861 38945 32864
rect 38979 32892 38991 32895
rect 39482 32892 39488 32904
rect 38979 32864 39488 32892
rect 38979 32861 38991 32864
rect 38933 32855 38991 32861
rect 39482 32852 39488 32864
rect 39540 32852 39546 32904
rect 42334 32852 42340 32904
rect 42392 32892 42398 32904
rect 42702 32892 42708 32904
rect 42392 32864 42708 32892
rect 42392 32852 42398 32864
rect 42702 32852 42708 32864
rect 42760 32892 42766 32904
rect 42996 32901 43024 32932
rect 44634 32920 44640 32972
rect 44692 32960 44698 32972
rect 46198 32960 46204 32972
rect 44692 32932 45600 32960
rect 46159 32932 46204 32960
rect 44692 32920 44698 32932
rect 42797 32895 42855 32901
rect 42797 32892 42809 32895
rect 42760 32864 42809 32892
rect 42760 32852 42766 32864
rect 42797 32861 42809 32864
rect 42843 32861 42855 32895
rect 42797 32855 42855 32861
rect 42981 32895 43039 32901
rect 42981 32861 42993 32895
rect 43027 32861 43039 32895
rect 43199 32895 43257 32901
rect 42981 32855 43039 32861
rect 43074 32873 43132 32879
rect 37274 32824 37280 32836
rect 35667 32796 35848 32824
rect 36004 32796 37280 32824
rect 35667 32793 35679 32796
rect 35621 32787 35679 32793
rect 29638 32716 29644 32768
rect 29696 32756 29702 32768
rect 29825 32759 29883 32765
rect 29825 32756 29837 32759
rect 29696 32728 29837 32756
rect 29696 32716 29702 32728
rect 29825 32725 29837 32728
rect 29871 32725 29883 32759
rect 35820 32756 35848 32796
rect 37274 32784 37280 32796
rect 37332 32784 37338 32836
rect 37553 32827 37611 32833
rect 37553 32793 37565 32827
rect 37599 32824 37611 32827
rect 37642 32824 37648 32836
rect 37599 32796 37648 32824
rect 37599 32793 37611 32796
rect 37553 32787 37611 32793
rect 37642 32784 37648 32796
rect 37700 32824 37706 32836
rect 40402 32824 40408 32836
rect 37700 32796 38792 32824
rect 40363 32796 40408 32824
rect 37700 32784 37706 32796
rect 35986 32756 35992 32768
rect 35820 32728 35992 32756
rect 29825 32719 29883 32725
rect 35986 32716 35992 32728
rect 36044 32756 36050 32768
rect 38289 32759 38347 32765
rect 38289 32756 38301 32759
rect 36044 32728 38301 32756
rect 36044 32716 36050 32728
rect 38289 32725 38301 32728
rect 38335 32756 38347 32759
rect 38654 32756 38660 32768
rect 38335 32728 38660 32756
rect 38335 32725 38347 32728
rect 38289 32719 38347 32725
rect 38654 32716 38660 32728
rect 38712 32716 38718 32768
rect 38764 32756 38792 32796
rect 40402 32784 40408 32796
rect 40460 32784 40466 32836
rect 41414 32784 41420 32836
rect 41472 32784 41478 32836
rect 40586 32756 40592 32768
rect 38764 32728 40592 32756
rect 40586 32716 40592 32728
rect 40644 32716 40650 32768
rect 42794 32716 42800 32768
rect 42852 32756 42858 32768
rect 42996 32756 43024 32855
rect 43074 32839 43086 32873
rect 43120 32839 43132 32873
rect 43199 32861 43211 32895
rect 43245 32892 43257 32895
rect 43346 32892 43352 32904
rect 43245 32864 43352 32892
rect 43245 32861 43257 32864
rect 43199 32855 43257 32861
rect 43346 32852 43352 32864
rect 43404 32852 43410 32904
rect 44082 32852 44088 32904
rect 44140 32892 44146 32904
rect 44361 32895 44419 32901
rect 44361 32892 44373 32895
rect 44140 32864 44373 32892
rect 44140 32852 44146 32864
rect 44361 32861 44373 32864
rect 44407 32861 44419 32895
rect 44361 32855 44419 32861
rect 45189 32895 45247 32901
rect 45189 32861 45201 32895
rect 45235 32861 45247 32895
rect 45572 32892 45600 32932
rect 46198 32920 46204 32932
rect 46256 32920 46262 32972
rect 47320 32969 47348 33000
rect 48774 32988 48780 33040
rect 48832 33028 48838 33040
rect 48832 33000 49096 33028
rect 48832 32988 48838 33000
rect 47305 32963 47363 32969
rect 47305 32929 47317 32963
rect 47351 32929 47363 32963
rect 47305 32923 47363 32929
rect 47578 32920 47584 32972
rect 47636 32960 47642 32972
rect 48961 32963 49019 32969
rect 48961 32960 48973 32963
rect 47636 32932 48973 32960
rect 47636 32920 47642 32932
rect 48961 32929 48973 32932
rect 49007 32929 49019 32963
rect 48961 32923 49019 32929
rect 46293 32895 46351 32901
rect 46293 32892 46305 32895
rect 45572 32864 46305 32892
rect 45189 32855 45247 32861
rect 46293 32861 46305 32864
rect 46339 32892 46351 32895
rect 46842 32892 46848 32904
rect 46339 32864 46848 32892
rect 46339 32861 46351 32864
rect 46293 32855 46351 32861
rect 43074 32836 43132 32839
rect 43070 32784 43076 32836
rect 43128 32784 43134 32836
rect 43441 32827 43499 32833
rect 43441 32793 43453 32827
rect 43487 32824 43499 32827
rect 43530 32824 43536 32836
rect 43487 32796 43536 32824
rect 43487 32793 43499 32796
rect 43441 32787 43499 32793
rect 43530 32784 43536 32796
rect 43588 32824 43594 32836
rect 45204 32824 45232 32855
rect 46842 32852 46848 32864
rect 46900 32852 46906 32904
rect 47394 32892 47400 32904
rect 47355 32864 47400 32892
rect 47394 32852 47400 32864
rect 47452 32852 47458 32904
rect 48590 32852 48596 32904
rect 48648 32892 48654 32904
rect 48685 32895 48743 32901
rect 48685 32892 48697 32895
rect 48648 32864 48697 32892
rect 48648 32852 48654 32864
rect 48685 32861 48697 32864
rect 48731 32861 48743 32895
rect 48685 32855 48743 32861
rect 48777 32895 48835 32901
rect 48777 32861 48789 32895
rect 48823 32861 48835 32895
rect 48777 32855 48835 32861
rect 48406 32824 48412 32836
rect 43588 32796 48412 32824
rect 43588 32784 43594 32796
rect 48406 32784 48412 32796
rect 48464 32784 48470 32836
rect 48792 32824 48820 32855
rect 48608 32796 48820 32824
rect 48976 32824 49004 32923
rect 49068 32901 49096 33000
rect 50709 32963 50767 32969
rect 50709 32960 50721 32963
rect 49620 32932 50721 32960
rect 49620 32904 49648 32932
rect 50709 32929 50721 32932
rect 50755 32960 50767 32963
rect 51074 32960 51080 32972
rect 50755 32932 51080 32960
rect 50755 32929 50767 32932
rect 50709 32923 50767 32929
rect 51074 32920 51080 32932
rect 51132 32920 51138 32972
rect 49053 32895 49111 32901
rect 49053 32861 49065 32895
rect 49099 32861 49111 32895
rect 49602 32892 49608 32904
rect 49563 32864 49608 32892
rect 49053 32855 49111 32861
rect 49602 32852 49608 32864
rect 49660 32852 49666 32904
rect 49786 32892 49792 32904
rect 49747 32864 49792 32892
rect 49786 32852 49792 32864
rect 49844 32892 49850 32904
rect 51276 32901 51304 33068
rect 52273 33065 52285 33099
rect 52319 33096 52331 33099
rect 52362 33096 52368 33108
rect 52319 33068 52368 33096
rect 52319 33065 52331 33068
rect 52273 33059 52331 33065
rect 52362 33056 52368 33068
rect 52420 33056 52426 33108
rect 54481 33099 54539 33105
rect 54481 33065 54493 33099
rect 54527 33096 54539 33099
rect 54570 33096 54576 33108
rect 54527 33068 54576 33096
rect 54527 33065 54539 33068
rect 54481 33059 54539 33065
rect 54570 33056 54576 33068
rect 54628 33056 54634 33108
rect 55493 33099 55551 33105
rect 55493 33065 55505 33099
rect 55539 33096 55551 33099
rect 55582 33096 55588 33108
rect 55539 33068 55588 33096
rect 55539 33065 55551 33068
rect 55493 33059 55551 33065
rect 55582 33056 55588 33068
rect 55640 33056 55646 33108
rect 56597 33099 56655 33105
rect 56597 33065 56609 33099
rect 56643 33096 56655 33099
rect 56686 33096 56692 33108
rect 56643 33068 56692 33096
rect 56643 33065 56655 33068
rect 56597 33059 56655 33065
rect 55766 32988 55772 33040
rect 55824 33028 55830 33040
rect 56612 33028 56640 33059
rect 56686 33056 56692 33068
rect 56744 33056 56750 33108
rect 57514 33096 57520 33108
rect 57475 33068 57520 33096
rect 57514 33056 57520 33068
rect 57572 33096 57578 33108
rect 58253 33099 58311 33105
rect 58253 33096 58265 33099
rect 57572 33068 58265 33096
rect 57572 33056 57578 33068
rect 58253 33065 58265 33068
rect 58299 33065 58311 33099
rect 58253 33059 58311 33065
rect 55824 33000 56640 33028
rect 55824 32988 55830 33000
rect 52270 32920 52276 32972
rect 52328 32960 52334 32972
rect 56778 32960 56784 32972
rect 52328 32932 56784 32960
rect 52328 32920 52334 32932
rect 50525 32895 50583 32901
rect 50525 32892 50537 32895
rect 49844 32864 50537 32892
rect 49844 32852 49850 32864
rect 50525 32861 50537 32864
rect 50571 32861 50583 32895
rect 50525 32855 50583 32861
rect 51261 32895 51319 32901
rect 51261 32861 51273 32895
rect 51307 32892 51319 32895
rect 51721 32895 51779 32901
rect 51721 32892 51733 32895
rect 51307 32864 51733 32892
rect 51307 32861 51319 32864
rect 51261 32855 51319 32861
rect 51721 32861 51733 32864
rect 51767 32861 51779 32895
rect 51721 32855 51779 32861
rect 52457 32895 52515 32901
rect 52457 32861 52469 32895
rect 52503 32861 52515 32895
rect 52457 32855 52515 32861
rect 50706 32824 50712 32836
rect 48976 32796 50712 32824
rect 48608 32768 48636 32796
rect 50706 32784 50712 32796
rect 50764 32784 50770 32836
rect 51626 32784 51632 32836
rect 51684 32824 51690 32836
rect 52472 32824 52500 32855
rect 52546 32852 52552 32904
rect 52604 32892 52610 32904
rect 52748 32901 52776 32932
rect 52733 32895 52791 32901
rect 52604 32864 52649 32892
rect 52604 32852 52610 32864
rect 52733 32861 52745 32895
rect 52779 32861 52791 32895
rect 52733 32855 52791 32861
rect 52825 32895 52883 32901
rect 52825 32861 52837 32895
rect 52871 32892 52883 32895
rect 52914 32892 52920 32904
rect 52871 32864 52920 32892
rect 52871 32861 52883 32864
rect 52825 32855 52883 32861
rect 52914 32852 52920 32864
rect 52972 32852 52978 32904
rect 53926 32892 53932 32904
rect 53887 32864 53932 32892
rect 53926 32852 53932 32864
rect 53984 32852 53990 32904
rect 54036 32901 54064 32932
rect 54021 32895 54079 32901
rect 54021 32861 54033 32895
rect 54067 32861 54079 32895
rect 54021 32855 54079 32861
rect 54110 32852 54116 32904
rect 54168 32892 54174 32904
rect 54205 32895 54263 32901
rect 54205 32892 54217 32895
rect 54168 32864 54217 32892
rect 54168 32852 54174 32864
rect 54205 32861 54217 32864
rect 54251 32861 54263 32895
rect 54205 32855 54263 32861
rect 54294 32852 54300 32904
rect 54352 32892 54358 32904
rect 55677 32895 55735 32901
rect 54352 32864 54397 32892
rect 54352 32852 54358 32864
rect 55677 32861 55689 32895
rect 55723 32861 55735 32895
rect 55677 32855 55735 32861
rect 53558 32824 53564 32836
rect 51684 32796 53564 32824
rect 51684 32784 51690 32796
rect 53558 32784 53564 32796
rect 53616 32824 53622 32836
rect 55692 32824 55720 32855
rect 55766 32852 55772 32904
rect 55824 32892 55830 32904
rect 55968 32901 55996 32932
rect 56778 32920 56784 32932
rect 56836 32920 56842 32972
rect 57146 32960 57152 32972
rect 57107 32932 57152 32960
rect 57146 32920 57152 32932
rect 57204 32920 57210 32972
rect 57974 32920 57980 32972
rect 58032 32960 58038 32972
rect 58069 32963 58127 32969
rect 58069 32960 58081 32963
rect 58032 32932 58081 32960
rect 58032 32920 58038 32932
rect 58069 32929 58081 32932
rect 58115 32929 58127 32963
rect 58069 32923 58127 32929
rect 55953 32895 56011 32901
rect 55824 32864 55869 32892
rect 55824 32852 55830 32864
rect 55953 32861 55965 32895
rect 55999 32861 56011 32895
rect 55953 32855 56011 32861
rect 56045 32895 56103 32901
rect 56045 32861 56057 32895
rect 56091 32892 56103 32895
rect 56226 32892 56232 32904
rect 56091 32864 56232 32892
rect 56091 32861 56103 32864
rect 56045 32855 56103 32861
rect 56226 32852 56232 32864
rect 56284 32852 56290 32904
rect 57241 32895 57299 32901
rect 57241 32861 57253 32895
rect 57287 32861 57299 32895
rect 57241 32855 57299 32861
rect 57054 32824 57060 32836
rect 53616 32796 57060 32824
rect 53616 32784 53622 32796
rect 57054 32784 57060 32796
rect 57112 32784 57118 32836
rect 57256 32824 57284 32855
rect 57422 32852 57428 32904
rect 57480 32892 57486 32904
rect 58345 32895 58403 32901
rect 58345 32892 58357 32895
rect 57480 32864 58357 32892
rect 57480 32852 57486 32864
rect 58345 32861 58357 32864
rect 58391 32861 58403 32895
rect 58345 32855 58403 32861
rect 58250 32824 58256 32836
rect 57256 32796 58256 32824
rect 58250 32784 58256 32796
rect 58308 32784 58314 32836
rect 44450 32756 44456 32768
rect 42852 32728 43024 32756
rect 44411 32728 44456 32756
rect 42852 32716 42858 32728
rect 44450 32716 44456 32728
rect 44508 32716 44514 32768
rect 45278 32756 45284 32768
rect 45239 32728 45284 32756
rect 45278 32716 45284 32728
rect 45336 32716 45342 32768
rect 47765 32759 47823 32765
rect 47765 32725 47777 32759
rect 47811 32756 47823 32759
rect 47946 32756 47952 32768
rect 47811 32728 47952 32756
rect 47811 32725 47823 32728
rect 47765 32719 47823 32725
rect 47946 32716 47952 32728
rect 48004 32716 48010 32768
rect 48590 32716 48596 32768
rect 48648 32716 48654 32768
rect 52730 32716 52736 32768
rect 52788 32756 52794 32768
rect 53285 32759 53343 32765
rect 53285 32756 53297 32759
rect 52788 32728 53297 32756
rect 52788 32716 52794 32728
rect 53285 32725 53297 32728
rect 53331 32725 53343 32759
rect 53285 32719 53343 32725
rect 58069 32759 58127 32765
rect 58069 32725 58081 32759
rect 58115 32756 58127 32759
rect 58158 32756 58164 32768
rect 58115 32728 58164 32756
rect 58115 32725 58127 32728
rect 58069 32719 58127 32725
rect 58158 32716 58164 32728
rect 58216 32716 58222 32768
rect 1104 32666 58880 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 58880 32666
rect 1104 32592 58880 32614
rect 29730 32512 29736 32564
rect 29788 32512 29794 32564
rect 30282 32512 30288 32564
rect 30340 32552 30346 32564
rect 30929 32555 30987 32561
rect 30340 32524 30512 32552
rect 30340 32512 30346 32524
rect 28350 32484 28356 32496
rect 28311 32456 28356 32484
rect 28350 32444 28356 32456
rect 28408 32444 28414 32496
rect 29638 32444 29644 32496
rect 29696 32444 29702 32496
rect 29748 32484 29776 32512
rect 30190 32484 30196 32496
rect 29748 32456 30196 32484
rect 30190 32444 30196 32456
rect 30248 32484 30254 32496
rect 30248 32456 30420 32484
rect 30248 32444 30254 32456
rect 30392 32425 30420 32456
rect 30377 32419 30435 32425
rect 30377 32385 30389 32419
rect 30423 32385 30435 32419
rect 30484 32416 30512 32524
rect 30929 32521 30941 32555
rect 30975 32552 30987 32555
rect 31018 32552 31024 32564
rect 30975 32524 31024 32552
rect 30975 32521 30987 32524
rect 30929 32515 30987 32521
rect 31018 32512 31024 32524
rect 31076 32512 31082 32564
rect 31570 32512 31576 32564
rect 31628 32552 31634 32564
rect 32309 32555 32367 32561
rect 32309 32552 32321 32555
rect 31628 32524 32321 32552
rect 31628 32512 31634 32524
rect 32309 32521 32321 32524
rect 32355 32521 32367 32555
rect 32309 32515 32367 32521
rect 32858 32512 32864 32564
rect 32916 32552 32922 32564
rect 34698 32552 34704 32564
rect 32916 32524 34560 32552
rect 34659 32524 34704 32552
rect 32916 32512 32922 32524
rect 34238 32444 34244 32496
rect 34296 32444 34302 32496
rect 34532 32484 34560 32524
rect 34698 32512 34704 32524
rect 34756 32512 34762 32564
rect 35713 32555 35771 32561
rect 35713 32521 35725 32555
rect 35759 32552 35771 32555
rect 35802 32552 35808 32564
rect 35759 32524 35808 32552
rect 35759 32521 35771 32524
rect 35713 32515 35771 32521
rect 35802 32512 35808 32524
rect 35860 32552 35866 32564
rect 36078 32552 36084 32564
rect 35860 32524 36084 32552
rect 35860 32512 35866 32524
rect 36078 32512 36084 32524
rect 36136 32512 36142 32564
rect 37366 32552 37372 32564
rect 36464 32524 37372 32552
rect 34532 32456 36400 32484
rect 31021 32419 31079 32425
rect 31021 32416 31033 32419
rect 30484 32388 31033 32416
rect 30377 32379 30435 32385
rect 31021 32385 31033 32388
rect 31067 32416 31079 32419
rect 31481 32419 31539 32425
rect 31481 32416 31493 32419
rect 31067 32388 31493 32416
rect 31067 32385 31079 32388
rect 31021 32379 31079 32385
rect 31481 32385 31493 32388
rect 31527 32385 31539 32419
rect 31481 32379 31539 32385
rect 32493 32419 32551 32425
rect 32493 32385 32505 32419
rect 32539 32385 32551 32419
rect 32493 32379 32551 32385
rect 30101 32351 30159 32357
rect 30101 32317 30113 32351
rect 30147 32348 30159 32351
rect 32306 32348 32312 32360
rect 30147 32320 32312 32348
rect 30147 32317 30159 32320
rect 30101 32311 30159 32317
rect 32306 32308 32312 32320
rect 32364 32308 32370 32360
rect 32508 32212 32536 32379
rect 34882 32376 34888 32428
rect 34940 32416 34946 32428
rect 35437 32419 35495 32425
rect 35437 32416 35449 32419
rect 34940 32388 35449 32416
rect 34940 32376 34946 32388
rect 35437 32385 35449 32388
rect 35483 32416 35495 32419
rect 35526 32416 35532 32428
rect 35483 32388 35532 32416
rect 35483 32385 35495 32388
rect 35437 32379 35495 32385
rect 35526 32376 35532 32388
rect 35584 32376 35590 32428
rect 32950 32348 32956 32360
rect 32911 32320 32956 32348
rect 32950 32308 32956 32320
rect 33008 32308 33014 32360
rect 33229 32351 33287 32357
rect 33229 32317 33241 32351
rect 33275 32348 33287 32351
rect 36265 32351 36323 32357
rect 36265 32348 36277 32351
rect 33275 32320 36277 32348
rect 33275 32317 33287 32320
rect 33229 32311 33287 32317
rect 36265 32317 36277 32320
rect 36311 32317 36323 32351
rect 36372 32348 36400 32456
rect 36464 32425 36492 32524
rect 37366 32512 37372 32524
rect 37424 32512 37430 32564
rect 37550 32552 37556 32564
rect 37511 32524 37556 32552
rect 37550 32512 37556 32524
rect 37608 32512 37614 32564
rect 38013 32555 38071 32561
rect 38013 32521 38025 32555
rect 38059 32552 38071 32555
rect 38194 32552 38200 32564
rect 38059 32524 38200 32552
rect 38059 32521 38071 32524
rect 38013 32515 38071 32521
rect 38194 32512 38200 32524
rect 38252 32512 38258 32564
rect 38608 32512 38614 32564
rect 38666 32552 38672 32564
rect 39114 32552 39120 32564
rect 38666 32524 38976 32552
rect 39075 32524 39120 32552
rect 38666 32512 38672 32524
rect 36541 32487 36599 32493
rect 36541 32453 36553 32487
rect 36587 32484 36599 32487
rect 37274 32484 37280 32496
rect 36587 32456 37280 32484
rect 36587 32453 36599 32456
rect 36541 32447 36599 32453
rect 37274 32444 37280 32456
rect 37332 32444 37338 32496
rect 37384 32484 37412 32512
rect 37918 32484 37924 32496
rect 37384 32456 37924 32484
rect 37918 32444 37924 32456
rect 37976 32484 37982 32496
rect 38290 32487 38348 32493
rect 38290 32484 38302 32487
rect 37976 32456 38302 32484
rect 37976 32444 37982 32456
rect 38290 32453 38302 32456
rect 38336 32453 38348 32487
rect 38290 32447 38348 32453
rect 38381 32487 38439 32493
rect 38381 32453 38393 32487
rect 38427 32484 38439 32487
rect 38838 32484 38844 32496
rect 38427 32456 38844 32484
rect 38427 32453 38439 32456
rect 38381 32447 38439 32453
rect 38838 32444 38844 32456
rect 38896 32444 38902 32496
rect 38948 32484 38976 32524
rect 39114 32512 39120 32524
rect 39172 32512 39178 32564
rect 40402 32512 40408 32564
rect 40460 32552 40466 32564
rect 40773 32555 40831 32561
rect 40773 32552 40785 32555
rect 40460 32524 40785 32552
rect 40460 32512 40466 32524
rect 40773 32521 40785 32524
rect 40819 32521 40831 32555
rect 41598 32552 41604 32564
rect 40773 32515 40831 32521
rect 41386 32524 41604 32552
rect 39393 32487 39451 32493
rect 39393 32484 39405 32487
rect 38948 32456 39405 32484
rect 39393 32453 39405 32456
rect 39439 32484 39451 32487
rect 40497 32487 40555 32493
rect 39439 32456 40264 32484
rect 39439 32453 39451 32456
rect 39393 32447 39451 32453
rect 36449 32419 36507 32425
rect 36449 32385 36461 32419
rect 36495 32416 36507 32419
rect 36633 32419 36691 32425
rect 36495 32388 36584 32416
rect 36495 32385 36507 32388
rect 36449 32379 36507 32385
rect 36556 32360 36584 32388
rect 36633 32385 36645 32419
rect 36679 32385 36691 32419
rect 36633 32379 36691 32385
rect 36771 32419 36829 32425
rect 36771 32385 36783 32419
rect 36817 32416 36829 32419
rect 38198 32419 38256 32425
rect 36817 32388 37780 32416
rect 36817 32385 36829 32388
rect 36771 32379 36829 32385
rect 36372 32320 36492 32348
rect 36265 32311 36323 32317
rect 36464 32292 36492 32320
rect 36538 32308 36544 32360
rect 36596 32308 36602 32360
rect 36446 32240 36452 32292
rect 36504 32240 36510 32292
rect 36648 32280 36676 32379
rect 36906 32348 36912 32360
rect 36867 32320 36912 32348
rect 36906 32308 36912 32320
rect 36964 32308 36970 32360
rect 37752 32280 37780 32388
rect 38198 32385 38210 32419
rect 38244 32414 38256 32419
rect 38244 32386 38424 32414
rect 38244 32385 38256 32386
rect 38198 32379 38256 32385
rect 38396 32348 38424 32386
rect 38470 32376 38476 32428
rect 38528 32425 38534 32428
rect 38528 32419 38557 32425
rect 38545 32385 38557 32419
rect 38528 32379 38557 32385
rect 38528 32376 38534 32379
rect 38654 32376 38660 32428
rect 38712 32416 38718 32428
rect 39298 32416 39304 32428
rect 38712 32388 38757 32416
rect 38948 32406 39304 32416
rect 38840 32388 39304 32406
rect 38712 32376 38718 32388
rect 38840 32378 38976 32388
rect 38840 32348 38868 32378
rect 39298 32376 39304 32388
rect 39356 32376 39362 32428
rect 39485 32419 39543 32425
rect 39485 32385 39497 32419
rect 39531 32385 39543 32419
rect 39485 32379 39543 32385
rect 38396 32320 38868 32348
rect 39206 32308 39212 32360
rect 39264 32348 39270 32360
rect 39500 32348 39528 32379
rect 39574 32376 39580 32428
rect 39632 32425 39638 32428
rect 40236 32425 40264 32456
rect 40497 32453 40509 32487
rect 40543 32484 40555 32487
rect 41386 32484 41414 32524
rect 41598 32512 41604 32524
rect 41656 32512 41662 32564
rect 41785 32555 41843 32561
rect 41785 32521 41797 32555
rect 41831 32521 41843 32555
rect 41785 32515 41843 32521
rect 40543 32456 41414 32484
rect 41509 32487 41567 32493
rect 40543 32453 40555 32456
rect 40497 32447 40555 32453
rect 41509 32453 41521 32487
rect 41555 32484 41567 32487
rect 41800 32484 41828 32515
rect 42886 32512 42892 32564
rect 42944 32552 42950 32564
rect 43165 32555 43223 32561
rect 43165 32552 43177 32555
rect 42944 32524 43177 32552
rect 42944 32512 42950 32524
rect 43165 32521 43177 32524
rect 43211 32521 43223 32555
rect 43165 32515 43223 32521
rect 43714 32512 43720 32564
rect 43772 32552 43778 32564
rect 46017 32555 46075 32561
rect 46017 32552 46029 32555
rect 43772 32524 46029 32552
rect 43772 32512 43778 32524
rect 46017 32521 46029 32524
rect 46063 32552 46075 32555
rect 46569 32555 46627 32561
rect 46569 32552 46581 32555
rect 46063 32524 46581 32552
rect 46063 32521 46075 32524
rect 46017 32515 46075 32521
rect 46569 32521 46581 32524
rect 46615 32552 46627 32555
rect 46934 32552 46940 32564
rect 46615 32524 46940 32552
rect 46615 32521 46627 32524
rect 46569 32515 46627 32521
rect 46934 32512 46940 32524
rect 46992 32512 46998 32564
rect 47210 32552 47216 32564
rect 47171 32524 47216 32552
rect 47210 32512 47216 32524
rect 47268 32512 47274 32564
rect 49697 32555 49755 32561
rect 49697 32521 49709 32555
rect 49743 32552 49755 32555
rect 49786 32552 49792 32564
rect 49743 32524 49792 32552
rect 49743 32521 49755 32524
rect 49697 32515 49755 32521
rect 49786 32512 49792 32524
rect 49844 32512 49850 32564
rect 50798 32512 50804 32564
rect 50856 32552 50862 32564
rect 50856 32524 51074 32552
rect 50856 32512 50862 32524
rect 43993 32487 44051 32493
rect 43993 32484 44005 32487
rect 41555 32456 41736 32484
rect 41800 32456 44005 32484
rect 41555 32453 41567 32456
rect 41509 32447 41567 32453
rect 39632 32419 39661 32425
rect 39649 32385 39661 32419
rect 39632 32379 39661 32385
rect 40221 32419 40279 32425
rect 40221 32385 40233 32419
rect 40267 32385 40279 32419
rect 40402 32416 40408 32428
rect 40363 32388 40408 32416
rect 40221 32379 40279 32385
rect 39632 32376 39638 32379
rect 40402 32376 40408 32388
rect 40460 32376 40466 32428
rect 40586 32416 40592 32428
rect 40547 32388 40592 32416
rect 40586 32376 40592 32388
rect 40644 32376 40650 32428
rect 41233 32419 41291 32425
rect 41233 32385 41245 32419
rect 41279 32416 41291 32419
rect 41322 32416 41328 32428
rect 41279 32388 41328 32416
rect 41279 32385 41291 32388
rect 41233 32379 41291 32385
rect 41322 32376 41328 32388
rect 41380 32376 41386 32428
rect 41417 32419 41475 32425
rect 41417 32385 41429 32419
rect 41463 32385 41475 32419
rect 41417 32379 41475 32385
rect 41601 32419 41659 32425
rect 41601 32385 41613 32419
rect 41647 32385 41659 32419
rect 41601 32379 41659 32385
rect 39264 32320 39528 32348
rect 39761 32351 39819 32357
rect 39264 32308 39270 32320
rect 39761 32317 39773 32351
rect 39807 32317 39819 32351
rect 39761 32311 39819 32317
rect 39574 32280 39580 32292
rect 36648 32252 37688 32280
rect 37752 32252 39580 32280
rect 35342 32212 35348 32224
rect 32508 32184 35348 32212
rect 35342 32172 35348 32184
rect 35400 32172 35406 32224
rect 36262 32172 36268 32224
rect 36320 32212 36326 32224
rect 37550 32212 37556 32224
rect 36320 32184 37556 32212
rect 36320 32172 36326 32184
rect 37550 32172 37556 32184
rect 37608 32172 37614 32224
rect 37660 32212 37688 32252
rect 39574 32240 39580 32252
rect 39632 32240 39638 32292
rect 39776 32280 39804 32311
rect 39850 32308 39856 32360
rect 39908 32348 39914 32360
rect 41432 32348 41460 32379
rect 39908 32320 41460 32348
rect 39908 32308 39914 32320
rect 41230 32280 41236 32292
rect 39776 32252 41236 32280
rect 41230 32240 41236 32252
rect 41288 32240 41294 32292
rect 39206 32212 39212 32224
rect 37660 32184 39212 32212
rect 39206 32172 39212 32184
rect 39264 32172 39270 32224
rect 40218 32172 40224 32224
rect 40276 32212 40282 32224
rect 41616 32212 41644 32379
rect 41708 32348 41736 32456
rect 43993 32453 44005 32456
rect 44039 32453 44051 32487
rect 43993 32447 44051 32453
rect 44450 32444 44456 32496
rect 44508 32444 44514 32496
rect 45922 32484 45928 32496
rect 45388 32456 45928 32484
rect 42794 32416 42800 32428
rect 42755 32388 42800 32416
rect 42794 32376 42800 32388
rect 42852 32376 42858 32428
rect 42978 32416 42984 32428
rect 42939 32388 42984 32416
rect 42978 32376 42984 32388
rect 43036 32376 43042 32428
rect 43714 32416 43720 32428
rect 43675 32388 43720 32416
rect 43714 32376 43720 32388
rect 43772 32376 43778 32428
rect 45388 32348 45416 32456
rect 45922 32444 45928 32456
rect 45980 32444 45986 32496
rect 48406 32444 48412 32496
rect 48464 32484 48470 32496
rect 49418 32484 49424 32496
rect 48464 32456 49424 32484
rect 48464 32444 48470 32456
rect 46842 32376 46848 32428
rect 46900 32416 46906 32428
rect 48041 32419 48099 32425
rect 48041 32416 48053 32419
rect 46900 32388 48053 32416
rect 46900 32376 46906 32388
rect 48041 32385 48053 32388
rect 48087 32416 48099 32419
rect 48590 32416 48596 32428
rect 48087 32388 48596 32416
rect 48087 32385 48099 32388
rect 48041 32379 48099 32385
rect 48590 32376 48596 32388
rect 48648 32376 48654 32428
rect 49344 32425 49372 32456
rect 49418 32444 49424 32456
rect 49476 32444 49482 32496
rect 51046 32484 51074 32524
rect 51350 32512 51356 32564
rect 51408 32552 51414 32564
rect 51537 32555 51595 32561
rect 51537 32552 51549 32555
rect 51408 32524 51549 32552
rect 51408 32512 51414 32524
rect 51537 32521 51549 32524
rect 51583 32521 51595 32555
rect 51537 32515 51595 32521
rect 51994 32512 52000 32564
rect 52052 32552 52058 32564
rect 52730 32552 52736 32564
rect 52052 32524 52736 32552
rect 52052 32512 52058 32524
rect 52730 32512 52736 32524
rect 52788 32512 52794 32564
rect 52914 32552 52920 32564
rect 52875 32524 52920 32552
rect 52914 32512 52920 32524
rect 52972 32512 52978 32564
rect 53926 32512 53932 32564
rect 53984 32552 53990 32564
rect 54205 32555 54263 32561
rect 54205 32552 54217 32555
rect 53984 32524 54217 32552
rect 53984 32512 53990 32524
rect 54205 32521 54217 32524
rect 54251 32521 54263 32555
rect 56226 32552 56232 32564
rect 56187 32524 56232 32552
rect 54205 32515 54263 32521
rect 56226 32512 56232 32524
rect 56284 32512 56290 32564
rect 57146 32512 57152 32564
rect 57204 32552 57210 32564
rect 57241 32555 57299 32561
rect 57241 32552 57253 32555
rect 57204 32524 57253 32552
rect 57204 32512 57210 32524
rect 57241 32521 57253 32524
rect 57287 32521 57299 32555
rect 57241 32515 57299 32521
rect 51813 32487 51871 32493
rect 51813 32484 51825 32487
rect 51046 32456 51825 32484
rect 51813 32453 51825 32456
rect 51859 32453 51871 32487
rect 51813 32447 51871 32453
rect 52564 32456 53236 32484
rect 49329 32419 49387 32425
rect 49329 32385 49341 32419
rect 49375 32385 49387 32419
rect 50706 32416 50712 32428
rect 50667 32388 50712 32416
rect 49329 32379 49387 32385
rect 50706 32376 50712 32388
rect 50764 32376 50770 32428
rect 50801 32419 50859 32425
rect 50801 32385 50813 32419
rect 50847 32385 50859 32419
rect 50801 32379 50859 32385
rect 41708 32320 45416 32348
rect 45465 32351 45523 32357
rect 45465 32317 45477 32351
rect 45511 32348 45523 32351
rect 46014 32348 46020 32360
rect 45511 32320 46020 32348
rect 45511 32317 45523 32320
rect 45465 32311 45523 32317
rect 46014 32308 46020 32320
rect 46072 32308 46078 32360
rect 47118 32308 47124 32360
rect 47176 32348 47182 32360
rect 47765 32351 47823 32357
rect 47765 32348 47777 32351
rect 47176 32320 47777 32348
rect 47176 32308 47182 32320
rect 47765 32317 47777 32320
rect 47811 32317 47823 32351
rect 47765 32311 47823 32317
rect 49421 32351 49479 32357
rect 49421 32317 49433 32351
rect 49467 32348 49479 32351
rect 50433 32351 50491 32357
rect 50433 32348 50445 32351
rect 49467 32320 50445 32348
rect 49467 32317 49479 32320
rect 49421 32311 49479 32317
rect 50433 32317 50445 32320
rect 50479 32317 50491 32351
rect 50816 32348 50844 32379
rect 50890 32376 50896 32428
rect 50948 32416 50954 32428
rect 50948 32388 50993 32416
rect 50948 32376 50954 32388
rect 51074 32376 51080 32428
rect 51132 32416 51138 32428
rect 51132 32388 51177 32416
rect 51132 32376 51138 32388
rect 51626 32376 51632 32428
rect 51684 32425 51690 32428
rect 51684 32419 51733 32425
rect 51684 32385 51687 32419
rect 51721 32385 51733 32419
rect 51902 32416 51908 32428
rect 51863 32388 51908 32416
rect 51684 32379 51733 32385
rect 51684 32376 51690 32379
rect 51902 32376 51908 32388
rect 51960 32376 51966 32428
rect 51994 32376 52000 32428
rect 52052 32425 52058 32428
rect 52052 32419 52091 32425
rect 52079 32385 52091 32419
rect 52052 32379 52091 32385
rect 52052 32376 52058 32379
rect 52178 32376 52184 32428
rect 52236 32416 52242 32428
rect 52236 32388 52281 32416
rect 52236 32376 52242 32388
rect 52564 32360 52592 32456
rect 52638 32376 52644 32428
rect 52696 32416 52702 32428
rect 53208 32425 53236 32456
rect 53374 32444 53380 32496
rect 53432 32484 53438 32496
rect 53561 32487 53619 32493
rect 53561 32484 53573 32487
rect 53432 32456 53573 32484
rect 53432 32444 53438 32456
rect 53561 32453 53573 32456
rect 53607 32453 53619 32487
rect 53561 32447 53619 32453
rect 54386 32444 54392 32496
rect 54444 32484 54450 32496
rect 54849 32487 54907 32493
rect 54849 32484 54861 32487
rect 54444 32456 54861 32484
rect 54444 32444 54450 32456
rect 54849 32453 54861 32456
rect 54895 32453 54907 32487
rect 54849 32447 54907 32453
rect 54938 32444 54944 32496
rect 54996 32484 55002 32496
rect 55677 32487 55735 32493
rect 55677 32484 55689 32487
rect 54996 32456 55689 32484
rect 54996 32444 55002 32456
rect 55677 32453 55689 32456
rect 55723 32453 55735 32487
rect 55677 32447 55735 32453
rect 55766 32444 55772 32496
rect 55824 32484 55830 32496
rect 55824 32456 56088 32484
rect 55824 32444 55830 32456
rect 53101 32419 53159 32425
rect 53101 32416 53113 32419
rect 52696 32388 53113 32416
rect 52696 32376 52702 32388
rect 53101 32385 53113 32388
rect 53147 32385 53159 32419
rect 53101 32379 53159 32385
rect 53193 32419 53251 32425
rect 53193 32385 53205 32419
rect 53239 32416 53251 32419
rect 53469 32419 53527 32425
rect 53239 32388 53420 32416
rect 53239 32385 53251 32388
rect 53193 32379 53251 32385
rect 50982 32348 50988 32360
rect 50816 32320 50988 32348
rect 50433 32311 50491 32317
rect 50982 32308 50988 32320
rect 51040 32308 51046 32360
rect 52546 32308 52552 32360
rect 52604 32308 52610 32360
rect 53116 32348 53144 32379
rect 53282 32348 53288 32360
rect 53116 32320 53288 32348
rect 53282 32308 53288 32320
rect 53340 32308 53346 32360
rect 47857 32283 47915 32289
rect 47857 32249 47869 32283
rect 47903 32280 47915 32283
rect 52270 32280 52276 32292
rect 47903 32252 52276 32280
rect 47903 32249 47915 32252
rect 47857 32243 47915 32249
rect 52270 32240 52276 32252
rect 52328 32240 52334 32292
rect 53392 32280 53420 32388
rect 53469 32385 53481 32419
rect 53515 32416 53527 32419
rect 53650 32416 53656 32428
rect 53515 32388 53656 32416
rect 53515 32385 53527 32388
rect 53469 32379 53527 32385
rect 53650 32376 53656 32388
rect 53708 32376 53714 32428
rect 54481 32419 54539 32425
rect 54481 32385 54493 32419
rect 54527 32416 54539 32419
rect 54570 32416 54576 32428
rect 54527 32388 54576 32416
rect 54527 32385 54539 32388
rect 54481 32379 54539 32385
rect 54570 32376 54576 32388
rect 54628 32376 54634 32428
rect 55582 32416 55588 32428
rect 55543 32388 55588 32416
rect 55582 32376 55588 32388
rect 55640 32376 55646 32428
rect 54110 32308 54116 32360
rect 54168 32348 54174 32360
rect 54389 32351 54447 32357
rect 54389 32348 54401 32351
rect 54168 32320 54401 32348
rect 54168 32308 54174 32320
rect 54389 32317 54401 32320
rect 54435 32317 54447 32351
rect 54389 32311 54447 32317
rect 54757 32351 54815 32357
rect 54757 32317 54769 32351
rect 54803 32348 54815 32351
rect 55784 32348 55812 32444
rect 55950 32416 55956 32428
rect 55911 32388 55956 32416
rect 55950 32376 55956 32388
rect 56008 32376 56014 32428
rect 56060 32425 56088 32456
rect 56318 32444 56324 32496
rect 56376 32484 56382 32496
rect 57330 32484 57336 32496
rect 56376 32456 57336 32484
rect 56376 32444 56382 32456
rect 56045 32419 56103 32425
rect 56045 32385 56057 32419
rect 56091 32385 56103 32419
rect 56045 32379 56103 32385
rect 56410 32376 56416 32428
rect 56468 32416 56474 32428
rect 56689 32419 56747 32425
rect 56689 32416 56701 32419
rect 56468 32388 56701 32416
rect 56468 32376 56474 32388
rect 56689 32385 56701 32388
rect 56735 32385 56747 32419
rect 56689 32379 56747 32385
rect 56778 32376 56784 32428
rect 56836 32416 56842 32428
rect 56980 32425 57008 32456
rect 57330 32444 57336 32456
rect 57388 32444 57394 32496
rect 56965 32419 57023 32425
rect 56836 32388 56881 32416
rect 56836 32376 56842 32388
rect 56965 32385 56977 32419
rect 57011 32385 57023 32419
rect 56965 32379 57023 32385
rect 57054 32376 57060 32428
rect 57112 32416 57118 32428
rect 57112 32388 57157 32416
rect 57112 32376 57118 32388
rect 54803 32320 55812 32348
rect 54803 32317 54815 32320
rect 54757 32311 54815 32317
rect 55950 32280 55956 32292
rect 53392 32252 55956 32280
rect 55950 32240 55956 32252
rect 56008 32240 56014 32292
rect 40276 32184 41644 32212
rect 40276 32172 40282 32184
rect 48130 32172 48136 32224
rect 48188 32212 48194 32224
rect 48225 32215 48283 32221
rect 48225 32212 48237 32215
rect 48188 32184 48237 32212
rect 48188 32172 48194 32184
rect 48225 32181 48237 32184
rect 48271 32181 48283 32215
rect 48225 32175 48283 32181
rect 49510 32172 49516 32224
rect 49568 32212 49574 32224
rect 52362 32212 52368 32224
rect 49568 32184 52368 32212
rect 49568 32172 49574 32184
rect 52362 32172 52368 32184
rect 52420 32172 52426 32224
rect 52638 32172 52644 32224
rect 52696 32212 52702 32224
rect 53650 32212 53656 32224
rect 52696 32184 53656 32212
rect 52696 32172 52702 32184
rect 53650 32172 53656 32184
rect 53708 32172 53714 32224
rect 57974 32172 57980 32224
rect 58032 32212 58038 32224
rect 58069 32215 58127 32221
rect 58069 32212 58081 32215
rect 58032 32184 58081 32212
rect 58032 32172 58038 32184
rect 58069 32181 58081 32184
rect 58115 32181 58127 32215
rect 58069 32175 58127 32181
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 30282 31968 30288 32020
rect 30340 32008 30346 32020
rect 30377 32011 30435 32017
rect 30377 32008 30389 32011
rect 30340 31980 30389 32008
rect 30340 31968 30346 31980
rect 30377 31977 30389 31980
rect 30423 31977 30435 32011
rect 30377 31971 30435 31977
rect 31110 31968 31116 32020
rect 31168 32008 31174 32020
rect 31205 32011 31263 32017
rect 31205 32008 31217 32011
rect 31168 31980 31217 32008
rect 31168 31968 31174 31980
rect 31205 31977 31217 31980
rect 31251 31977 31263 32011
rect 31205 31971 31263 31977
rect 32306 31968 32312 32020
rect 32364 32008 32370 32020
rect 34149 32011 34207 32017
rect 32364 31980 34100 32008
rect 32364 31968 32370 31980
rect 30190 31900 30196 31952
rect 30248 31940 30254 31952
rect 34072 31940 34100 31980
rect 34149 31977 34161 32011
rect 34195 32008 34207 32011
rect 34238 32008 34244 32020
rect 34195 31980 34244 32008
rect 34195 31977 34207 31980
rect 34149 31971 34207 31977
rect 34238 31968 34244 31980
rect 34296 31968 34302 32020
rect 35342 32008 35348 32020
rect 35303 31980 35348 32008
rect 35342 31968 35348 31980
rect 35400 31968 35406 32020
rect 36354 31968 36360 32020
rect 36412 32008 36418 32020
rect 36541 32011 36599 32017
rect 36541 32008 36553 32011
rect 36412 31980 36553 32008
rect 36412 31968 36418 31980
rect 36541 31977 36553 31980
rect 36587 31977 36599 32011
rect 36541 31971 36599 31977
rect 37274 31968 37280 32020
rect 37332 32008 37338 32020
rect 38470 32008 38476 32020
rect 37332 31980 38476 32008
rect 37332 31968 37338 31980
rect 38470 31968 38476 31980
rect 38528 31968 38534 32020
rect 38562 31968 38568 32020
rect 38620 32008 38626 32020
rect 38654 32008 38660 32020
rect 38620 31980 38660 32008
rect 38620 31968 38626 31980
rect 38654 31968 38660 31980
rect 38712 32008 38718 32020
rect 38749 32011 38807 32017
rect 38749 32008 38761 32011
rect 38712 31980 38761 32008
rect 38712 31968 38718 31980
rect 38749 31977 38761 31980
rect 38795 31977 38807 32011
rect 38749 31971 38807 31977
rect 41141 32011 41199 32017
rect 41141 31977 41153 32011
rect 41187 32008 41199 32011
rect 41230 32008 41236 32020
rect 41187 31980 41236 32008
rect 41187 31977 41199 31980
rect 41141 31971 41199 31977
rect 41230 31968 41236 31980
rect 41288 31968 41294 32020
rect 41598 32008 41604 32020
rect 41559 31980 41604 32008
rect 41598 31968 41604 31980
rect 41656 31968 41662 32020
rect 42886 31968 42892 32020
rect 42944 32008 42950 32020
rect 43898 32008 43904 32020
rect 42944 31980 43904 32008
rect 42944 31968 42950 31980
rect 43898 31968 43904 31980
rect 43956 31968 43962 32020
rect 46934 32008 46940 32020
rect 46895 31980 46940 32008
rect 46934 31968 46940 31980
rect 46992 32008 46998 32020
rect 47762 32008 47768 32020
rect 46992 31980 47768 32008
rect 46992 31968 46998 31980
rect 47762 31968 47768 31980
rect 47820 31968 47826 32020
rect 48130 32008 48136 32020
rect 48091 31980 48136 32008
rect 48130 31968 48136 31980
rect 48188 31968 48194 32020
rect 48682 31968 48688 32020
rect 48740 32008 48746 32020
rect 49050 32008 49056 32020
rect 48740 31980 49056 32008
rect 48740 31968 48746 31980
rect 49050 31968 49056 31980
rect 49108 32008 49114 32020
rect 49421 32011 49479 32017
rect 49421 32008 49433 32011
rect 49108 31980 49433 32008
rect 49108 31968 49114 31980
rect 49421 31977 49433 31980
rect 49467 31977 49479 32011
rect 49421 31971 49479 31977
rect 50985 32011 51043 32017
rect 50985 31977 50997 32011
rect 51031 32008 51043 32011
rect 52178 32008 52184 32020
rect 51031 31980 52184 32008
rect 51031 31977 51043 31980
rect 50985 31971 51043 31977
rect 52178 31968 52184 31980
rect 52236 31968 52242 32020
rect 53374 32008 53380 32020
rect 52380 31980 53380 32008
rect 40037 31943 40095 31949
rect 40037 31940 40049 31943
rect 30248 31912 31340 31940
rect 34072 31912 40049 31940
rect 30248 31900 30254 31912
rect 31312 31872 31340 31912
rect 40037 31909 40049 31912
rect 40083 31909 40095 31943
rect 40037 31903 40095 31909
rect 42426 31900 42432 31952
rect 42484 31940 42490 31952
rect 43625 31943 43683 31949
rect 43625 31940 43637 31943
rect 42484 31912 43637 31940
rect 42484 31900 42490 31912
rect 43625 31909 43637 31912
rect 43671 31909 43683 31943
rect 43625 31903 43683 31909
rect 47578 31900 47584 31952
rect 47636 31940 47642 31952
rect 47636 31912 48912 31940
rect 47636 31900 47642 31912
rect 32950 31872 32956 31884
rect 31312 31844 32956 31872
rect 32950 31832 32956 31844
rect 33008 31832 33014 31884
rect 33505 31875 33563 31881
rect 33505 31841 33517 31875
rect 33551 31872 33563 31875
rect 34606 31872 34612 31884
rect 33551 31844 34612 31872
rect 33551 31841 33563 31844
rect 33505 31835 33563 31841
rect 34606 31832 34612 31844
rect 34664 31832 34670 31884
rect 35342 31832 35348 31884
rect 35400 31872 35406 31884
rect 35526 31872 35532 31884
rect 35400 31844 35532 31872
rect 35400 31832 35406 31844
rect 35526 31832 35532 31844
rect 35584 31832 35590 31884
rect 35805 31875 35863 31881
rect 35805 31841 35817 31875
rect 35851 31872 35863 31875
rect 35894 31872 35900 31884
rect 35851 31844 35900 31872
rect 35851 31841 35863 31844
rect 35805 31835 35863 31841
rect 35894 31832 35900 31844
rect 35952 31832 35958 31884
rect 35989 31875 36047 31881
rect 35989 31841 36001 31875
rect 36035 31872 36047 31875
rect 36078 31872 36084 31884
rect 36035 31844 36084 31872
rect 36035 31841 36047 31844
rect 35989 31835 36047 31841
rect 36078 31832 36084 31844
rect 36136 31832 36142 31884
rect 36262 31832 36268 31884
rect 36320 31832 36326 31884
rect 37274 31872 37280 31884
rect 36832 31844 37280 31872
rect 29917 31807 29975 31813
rect 29917 31773 29929 31807
rect 29963 31804 29975 31807
rect 30282 31804 30288 31816
rect 29963 31776 30288 31804
rect 29963 31773 29975 31776
rect 29917 31767 29975 31773
rect 30282 31764 30288 31776
rect 30340 31764 30346 31816
rect 33597 31807 33655 31813
rect 33597 31773 33609 31807
rect 33643 31804 33655 31807
rect 34241 31807 34299 31813
rect 34241 31804 34253 31807
rect 33643 31776 34253 31804
rect 33643 31773 33655 31776
rect 33597 31767 33655 31773
rect 34241 31773 34253 31776
rect 34287 31804 34299 31807
rect 34698 31804 34704 31816
rect 34287 31776 34704 31804
rect 34287 31773 34299 31776
rect 34241 31767 34299 31773
rect 34698 31764 34704 31776
rect 34756 31764 34762 31816
rect 36280 31804 36308 31832
rect 35866 31776 36308 31804
rect 32398 31736 32404 31748
rect 32246 31708 32404 31736
rect 32398 31696 32404 31708
rect 32456 31696 32462 31748
rect 32674 31736 32680 31748
rect 32635 31708 32680 31736
rect 32674 31696 32680 31708
rect 32732 31696 32738 31748
rect 35713 31739 35771 31745
rect 35713 31705 35725 31739
rect 35759 31736 35771 31739
rect 35866 31736 35894 31776
rect 36538 31764 36544 31816
rect 36596 31804 36602 31816
rect 36722 31804 36728 31816
rect 36596 31776 36728 31804
rect 36596 31764 36602 31776
rect 36722 31764 36728 31776
rect 36780 31764 36786 31816
rect 36832 31813 36860 31844
rect 37274 31832 37280 31844
rect 37332 31832 37338 31884
rect 38286 31872 38292 31884
rect 37384 31844 38292 31872
rect 36817 31807 36875 31813
rect 36817 31773 36829 31807
rect 36863 31773 36875 31807
rect 37182 31804 37188 31816
rect 37143 31776 37188 31804
rect 36817 31767 36875 31773
rect 37182 31764 37188 31776
rect 37240 31764 37246 31816
rect 37384 31804 37412 31844
rect 38286 31832 38292 31844
rect 38344 31832 38350 31884
rect 42150 31872 42156 31884
rect 40512 31844 42156 31872
rect 37292 31776 37412 31804
rect 35759 31708 35894 31736
rect 36909 31739 36967 31745
rect 35759 31705 35771 31708
rect 35713 31699 35771 31705
rect 36909 31705 36921 31739
rect 36955 31705 36967 31739
rect 36909 31699 36967 31705
rect 37047 31739 37105 31745
rect 37047 31705 37059 31739
rect 37093 31736 37105 31739
rect 37292 31736 37320 31776
rect 37550 31764 37556 31816
rect 37608 31804 37614 31816
rect 37645 31807 37703 31813
rect 37645 31804 37657 31807
rect 37608 31776 37657 31804
rect 37608 31764 37614 31776
rect 37645 31773 37657 31776
rect 37691 31773 37703 31807
rect 40218 31804 40224 31816
rect 40179 31776 40224 31804
rect 37645 31767 37703 31773
rect 40218 31764 40224 31776
rect 40276 31764 40282 31816
rect 40402 31804 40408 31816
rect 40363 31776 40408 31804
rect 40402 31764 40408 31776
rect 40460 31764 40466 31816
rect 38838 31736 38844 31748
rect 37093 31708 37320 31736
rect 37384 31708 38844 31736
rect 37093 31705 37105 31708
rect 37047 31699 37105 31705
rect 29822 31668 29828 31680
rect 29783 31640 29828 31668
rect 29822 31628 29828 31640
rect 29880 31628 29886 31680
rect 35802 31628 35808 31680
rect 35860 31668 35866 31680
rect 36262 31668 36268 31680
rect 35860 31640 36268 31668
rect 35860 31628 35866 31640
rect 36262 31628 36268 31640
rect 36320 31628 36326 31680
rect 36814 31628 36820 31680
rect 36872 31668 36878 31680
rect 36924 31668 36952 31699
rect 37384 31668 37412 31708
rect 38838 31696 38844 31708
rect 38896 31736 38902 31748
rect 40034 31736 40040 31748
rect 38896 31708 40040 31736
rect 38896 31696 38902 31708
rect 40034 31696 40040 31708
rect 40092 31696 40098 31748
rect 40313 31739 40371 31745
rect 40313 31705 40325 31739
rect 40359 31736 40371 31739
rect 40512 31736 40540 31844
rect 42150 31832 42156 31844
rect 42208 31832 42214 31884
rect 42886 31832 42892 31884
rect 42944 31872 42950 31884
rect 43254 31872 43260 31884
rect 42944 31844 43260 31872
rect 42944 31832 42950 31844
rect 43254 31832 43260 31844
rect 43312 31832 43318 31884
rect 45833 31875 45891 31881
rect 45833 31841 45845 31875
rect 45879 31872 45891 31875
rect 47210 31872 47216 31884
rect 45879 31844 47216 31872
rect 45879 31841 45891 31844
rect 45833 31835 45891 31841
rect 47210 31832 47216 31844
rect 47268 31832 47274 31884
rect 47670 31832 47676 31884
rect 47728 31872 47734 31884
rect 47949 31875 48007 31881
rect 47949 31872 47961 31875
rect 47728 31844 47961 31872
rect 47728 31832 47734 31844
rect 47949 31841 47961 31844
rect 47995 31841 48007 31875
rect 48777 31875 48835 31881
rect 48777 31872 48789 31875
rect 47949 31835 48007 31841
rect 48240 31844 48789 31872
rect 48240 31816 48268 31844
rect 48777 31841 48789 31844
rect 48823 31841 48835 31875
rect 48777 31835 48835 31841
rect 40589 31807 40647 31813
rect 40589 31773 40601 31807
rect 40635 31804 40647 31807
rect 41322 31804 41328 31816
rect 40635 31776 41328 31804
rect 40635 31773 40647 31776
rect 40589 31767 40647 31773
rect 41322 31764 41328 31776
rect 41380 31764 41386 31816
rect 42794 31764 42800 31816
rect 42852 31804 42858 31816
rect 42981 31807 43039 31813
rect 42981 31804 42993 31807
rect 42852 31776 42993 31804
rect 42852 31764 42858 31776
rect 42981 31773 42993 31776
rect 43027 31773 43039 31807
rect 42981 31767 43039 31773
rect 43070 31764 43076 31816
rect 43128 31804 43134 31816
rect 43165 31807 43223 31813
rect 43165 31804 43177 31807
rect 43128 31776 43177 31804
rect 43128 31764 43134 31776
rect 43165 31773 43177 31776
rect 43211 31773 43223 31807
rect 44266 31804 44272 31816
rect 44227 31776 44272 31804
rect 43165 31767 43223 31773
rect 44266 31764 44272 31776
rect 44324 31764 44330 31816
rect 45922 31804 45928 31816
rect 45883 31776 45928 31804
rect 45922 31764 45928 31776
rect 45980 31764 45986 31816
rect 48222 31804 48228 31816
rect 48183 31776 48228 31804
rect 48222 31764 48228 31776
rect 48280 31764 48286 31816
rect 48590 31764 48596 31816
rect 48648 31804 48654 31816
rect 48884 31813 48912 31912
rect 51902 31900 51908 31952
rect 51960 31940 51966 31952
rect 52380 31940 52408 31980
rect 53374 31968 53380 31980
rect 53432 31968 53438 32020
rect 53745 32011 53803 32017
rect 53745 31977 53757 32011
rect 53791 32008 53803 32011
rect 54478 32008 54484 32020
rect 53791 31980 54484 32008
rect 53791 31977 53803 31980
rect 53745 31971 53803 31977
rect 54478 31968 54484 31980
rect 54536 31968 54542 32020
rect 56410 32008 56416 32020
rect 56371 31980 56416 32008
rect 56410 31968 56416 31980
rect 56468 31968 56474 32020
rect 51960 31912 52408 31940
rect 52457 31943 52515 31949
rect 51960 31900 51966 31912
rect 52457 31909 52469 31943
rect 52503 31940 52515 31943
rect 52503 31912 53144 31940
rect 52503 31909 52515 31912
rect 52457 31903 52515 31909
rect 50890 31872 50896 31884
rect 50724 31844 50896 31872
rect 50724 31813 50752 31844
rect 50890 31832 50896 31844
rect 50948 31872 50954 31884
rect 51537 31875 51595 31881
rect 52365 31880 52423 31881
rect 51537 31872 51549 31875
rect 50948 31844 51549 31872
rect 50948 31832 50954 31844
rect 51537 31841 51549 31844
rect 51583 31872 51595 31875
rect 52288 31875 52423 31880
rect 52288 31872 52377 31875
rect 51583 31852 52377 31872
rect 51583 31844 52316 31852
rect 51583 31841 51595 31844
rect 51537 31835 51595 31841
rect 52365 31841 52377 31852
rect 52411 31841 52423 31875
rect 52365 31835 52423 31841
rect 48685 31807 48743 31813
rect 48685 31804 48697 31807
rect 48648 31776 48697 31804
rect 48648 31764 48654 31776
rect 48685 31773 48697 31776
rect 48731 31804 48743 31807
rect 48869 31807 48927 31813
rect 48731 31776 48820 31804
rect 48731 31773 48743 31776
rect 48685 31767 48743 31773
rect 40359 31708 40540 31736
rect 40359 31705 40371 31708
rect 40313 31699 40371 31705
rect 42886 31696 42892 31748
rect 42944 31736 42950 31748
rect 42944 31708 44404 31736
rect 42944 31696 42950 31708
rect 36872 31640 37412 31668
rect 38289 31671 38347 31677
rect 36872 31628 36878 31640
rect 38289 31637 38301 31671
rect 38335 31668 38347 31671
rect 38930 31668 38936 31680
rect 38335 31640 38936 31668
rect 38335 31637 38347 31640
rect 38289 31631 38347 31637
rect 38930 31628 38936 31640
rect 38988 31628 38994 31680
rect 39022 31628 39028 31680
rect 39080 31668 39086 31680
rect 39301 31671 39359 31677
rect 39301 31668 39313 31671
rect 39080 31640 39313 31668
rect 39080 31628 39086 31640
rect 39301 31637 39313 31640
rect 39347 31637 39359 31671
rect 43070 31668 43076 31680
rect 43031 31640 43076 31668
rect 39301 31631 39359 31637
rect 43070 31628 43076 31640
rect 43128 31628 43134 31680
rect 44376 31677 44404 31708
rect 45554 31696 45560 31748
rect 45612 31736 45618 31748
rect 46014 31736 46020 31748
rect 45612 31708 46020 31736
rect 45612 31696 45618 31708
rect 46014 31696 46020 31708
rect 46072 31696 46078 31748
rect 47854 31736 47860 31748
rect 46216 31708 47860 31736
rect 44361 31671 44419 31677
rect 44361 31637 44373 31671
rect 44407 31637 44419 31671
rect 44361 31631 44419 31637
rect 45278 31628 45284 31680
rect 45336 31668 45342 31680
rect 46216 31668 46244 31708
rect 47854 31696 47860 31708
rect 47912 31696 47918 31748
rect 48792 31736 48820 31776
rect 48869 31773 48881 31807
rect 48915 31773 48927 31807
rect 49329 31807 49387 31813
rect 49329 31804 49341 31807
rect 48869 31767 48927 31773
rect 48976 31776 49341 31804
rect 48976 31736 49004 31776
rect 49329 31773 49341 31776
rect 49375 31773 49387 31807
rect 49329 31767 49387 31773
rect 50709 31807 50767 31813
rect 50709 31773 50721 31807
rect 50755 31773 50767 31807
rect 50982 31804 50988 31816
rect 50943 31776 50988 31804
rect 50709 31767 50767 31773
rect 50982 31764 50988 31776
rect 51040 31764 51046 31816
rect 51442 31804 51448 31816
rect 51403 31776 51448 31804
rect 51442 31764 51448 31776
rect 51500 31764 51506 31816
rect 51626 31804 51632 31816
rect 51587 31776 51632 31804
rect 51626 31764 51632 31776
rect 51684 31764 51690 31816
rect 52546 31804 52552 31816
rect 52288 31776 52552 31804
rect 50798 31736 50804 31748
rect 48792 31708 49004 31736
rect 50759 31708 50804 31736
rect 50798 31696 50804 31708
rect 50856 31696 50862 31748
rect 51000 31736 51028 31764
rect 52288 31736 52316 31776
rect 52546 31764 52552 31776
rect 52604 31764 52610 31816
rect 53116 31813 53144 31912
rect 53392 31872 53420 31968
rect 54570 31900 54576 31952
rect 54628 31940 54634 31952
rect 57885 31943 57943 31949
rect 54628 31912 57008 31940
rect 54628 31900 54634 31912
rect 54757 31875 54815 31881
rect 54757 31872 54769 31875
rect 53392 31844 54769 31872
rect 53282 31813 53288 31816
rect 52641 31807 52699 31813
rect 52641 31773 52653 31807
rect 52687 31773 52699 31807
rect 52641 31767 52699 31773
rect 53101 31807 53159 31813
rect 53101 31773 53113 31807
rect 53147 31773 53159 31807
rect 53101 31767 53159 31773
rect 53249 31807 53288 31813
rect 53249 31773 53261 31807
rect 53249 31767 53288 31773
rect 51000 31708 52316 31736
rect 52362 31696 52368 31748
rect 52420 31736 52426 31748
rect 52656 31736 52684 31767
rect 53282 31764 53288 31767
rect 53340 31764 53346 31816
rect 53392 31813 53420 31844
rect 54757 31841 54769 31844
rect 54803 31872 54815 31875
rect 54803 31844 55352 31872
rect 54803 31841 54815 31844
rect 54757 31835 54815 31841
rect 53377 31807 53435 31813
rect 53377 31773 53389 31807
rect 53423 31773 53435 31807
rect 53377 31767 53435 31773
rect 53558 31764 53564 31816
rect 53616 31813 53622 31816
rect 53616 31804 53624 31813
rect 54938 31804 54944 31816
rect 53616 31776 53661 31804
rect 54221 31776 54944 31804
rect 53616 31767 53624 31776
rect 53616 31764 53622 31767
rect 53469 31739 53527 31745
rect 53469 31736 53481 31739
rect 52420 31708 53481 31736
rect 52420 31696 52426 31708
rect 53469 31705 53481 31708
rect 53515 31736 53527 31739
rect 54221 31736 54249 31776
rect 54938 31764 54944 31776
rect 54996 31764 55002 31816
rect 55324 31804 55352 31844
rect 55398 31832 55404 31884
rect 55456 31872 55462 31884
rect 55861 31875 55919 31881
rect 55861 31872 55873 31875
rect 55456 31844 55873 31872
rect 55456 31832 55462 31844
rect 55861 31841 55873 31844
rect 55907 31841 55919 31875
rect 55861 31835 55919 31841
rect 56229 31875 56287 31881
rect 56229 31841 56241 31875
rect 56275 31872 56287 31875
rect 56318 31872 56324 31884
rect 56275 31844 56324 31872
rect 56275 31841 56287 31844
rect 56229 31835 56287 31841
rect 55582 31804 55588 31816
rect 55324 31776 55588 31804
rect 55582 31764 55588 31776
rect 55640 31804 55646 31816
rect 55769 31807 55827 31813
rect 55769 31804 55781 31807
rect 55640 31776 55781 31804
rect 55640 31764 55646 31776
rect 55769 31773 55781 31776
rect 55815 31773 55827 31807
rect 55769 31767 55827 31773
rect 53515 31708 54249 31736
rect 53515 31705 53527 31708
rect 53469 31699 53527 31705
rect 54386 31696 54392 31748
rect 54444 31736 54450 31748
rect 54573 31739 54631 31745
rect 54573 31736 54585 31739
rect 54444 31708 54585 31736
rect 54444 31696 54450 31708
rect 54573 31705 54585 31708
rect 54619 31705 54631 31739
rect 55876 31736 55904 31835
rect 56318 31832 56324 31844
rect 56376 31832 56382 31884
rect 55950 31764 55956 31816
rect 56008 31804 56014 31816
rect 56134 31804 56140 31816
rect 56008 31776 56140 31804
rect 56008 31764 56014 31776
rect 56134 31764 56140 31776
rect 56192 31804 56198 31816
rect 56873 31807 56931 31813
rect 56873 31804 56885 31807
rect 56192 31803 56364 31804
rect 56428 31803 56885 31804
rect 56192 31776 56885 31803
rect 56192 31764 56198 31776
rect 56336 31775 56456 31776
rect 56873 31773 56885 31776
rect 56919 31773 56931 31807
rect 56980 31804 57008 31912
rect 57885 31909 57897 31943
rect 57931 31940 57943 31943
rect 58066 31940 58072 31952
rect 57931 31912 58072 31940
rect 57931 31909 57943 31912
rect 57885 31903 57943 31909
rect 58066 31900 58072 31912
rect 58124 31900 58130 31952
rect 58342 31872 58348 31884
rect 57164 31844 58348 31872
rect 57057 31807 57115 31813
rect 57057 31804 57069 31807
rect 56980 31776 57069 31804
rect 56873 31767 56931 31773
rect 57057 31773 57069 31776
rect 57103 31773 57115 31807
rect 57057 31767 57115 31773
rect 57164 31736 57192 31844
rect 58342 31832 58348 31844
rect 58400 31832 58406 31884
rect 57606 31804 57612 31816
rect 57567 31776 57612 31804
rect 57606 31764 57612 31776
rect 57664 31764 57670 31816
rect 57701 31807 57759 31813
rect 57701 31773 57713 31807
rect 57747 31804 57759 31807
rect 58250 31804 58256 31816
rect 57747 31776 58256 31804
rect 57747 31773 57759 31776
rect 57701 31767 57759 31773
rect 58250 31764 58256 31776
rect 58308 31804 58314 31816
rect 58526 31804 58532 31816
rect 58308 31776 58532 31804
rect 58308 31764 58314 31776
rect 58526 31764 58532 31776
rect 58584 31764 58590 31816
rect 55876 31708 57192 31736
rect 54573 31699 54631 31705
rect 57790 31696 57796 31748
rect 57848 31736 57854 31748
rect 57885 31739 57943 31745
rect 57885 31736 57897 31739
rect 57848 31708 57897 31736
rect 57848 31696 57854 31708
rect 57885 31705 57897 31708
rect 57931 31705 57943 31739
rect 57885 31699 57943 31705
rect 46382 31668 46388 31680
rect 45336 31640 46244 31668
rect 46343 31640 46388 31668
rect 45336 31628 45342 31640
rect 46382 31628 46388 31640
rect 46440 31628 46446 31680
rect 47118 31628 47124 31680
rect 47176 31668 47182 31680
rect 47397 31671 47455 31677
rect 47397 31668 47409 31671
rect 47176 31640 47409 31668
rect 47176 31628 47182 31640
rect 47397 31637 47409 31640
rect 47443 31637 47455 31671
rect 47397 31631 47455 31637
rect 47578 31628 47584 31680
rect 47636 31668 47642 31680
rect 47949 31671 48007 31677
rect 47949 31668 47961 31671
rect 47636 31640 47961 31668
rect 47636 31628 47642 31640
rect 47949 31637 47961 31640
rect 47995 31637 48007 31671
rect 47949 31631 48007 31637
rect 55030 31628 55036 31680
rect 55088 31668 55094 31680
rect 57974 31668 57980 31680
rect 55088 31640 57980 31668
rect 55088 31628 55094 31640
rect 57974 31628 57980 31640
rect 58032 31628 58038 31680
rect 1104 31578 58880 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 58880 31578
rect 1104 31504 58880 31526
rect 28258 31424 28264 31476
rect 28316 31464 28322 31476
rect 28445 31467 28503 31473
rect 28445 31464 28457 31467
rect 28316 31436 28457 31464
rect 28316 31424 28322 31436
rect 28445 31433 28457 31436
rect 28491 31433 28503 31467
rect 32398 31464 32404 31476
rect 32359 31436 32404 31464
rect 28445 31427 28503 31433
rect 32398 31424 32404 31436
rect 32456 31424 32462 31476
rect 32674 31424 32680 31476
rect 32732 31464 32738 31476
rect 35069 31467 35127 31473
rect 32732 31436 35020 31464
rect 32732 31424 32738 31436
rect 29822 31396 29828 31408
rect 29486 31368 29828 31396
rect 29822 31356 29828 31368
rect 29880 31356 29886 31408
rect 29917 31399 29975 31405
rect 29917 31365 29929 31399
rect 29963 31396 29975 31399
rect 33870 31396 33876 31408
rect 29963 31368 33876 31396
rect 29963 31365 29975 31368
rect 29917 31359 29975 31365
rect 33870 31356 33876 31368
rect 33928 31356 33934 31408
rect 34606 31356 34612 31408
rect 34664 31356 34670 31408
rect 30190 31288 30196 31340
rect 30248 31328 30254 31340
rect 32493 31331 32551 31337
rect 30248 31300 30293 31328
rect 30248 31288 30254 31300
rect 32493 31297 32505 31331
rect 32539 31328 32551 31331
rect 32858 31328 32864 31340
rect 32539 31300 32864 31328
rect 32539 31297 32551 31300
rect 32493 31291 32551 31297
rect 32858 31288 32864 31300
rect 32916 31288 32922 31340
rect 32950 31288 32956 31340
rect 33008 31328 33014 31340
rect 33321 31331 33379 31337
rect 33321 31328 33333 31331
rect 33008 31300 33333 31328
rect 33008 31288 33014 31300
rect 33321 31297 33333 31300
rect 33367 31297 33379 31331
rect 34992 31328 35020 31436
rect 35069 31433 35081 31467
rect 35115 31464 35127 31467
rect 35342 31464 35348 31476
rect 35115 31436 35348 31464
rect 35115 31433 35127 31436
rect 35069 31427 35127 31433
rect 35342 31424 35348 31436
rect 35400 31424 35406 31476
rect 35897 31467 35955 31473
rect 35897 31433 35909 31467
rect 35943 31464 35955 31467
rect 36262 31464 36268 31476
rect 35943 31436 36268 31464
rect 35943 31433 35955 31436
rect 35897 31427 35955 31433
rect 36262 31424 36268 31436
rect 36320 31424 36326 31476
rect 38102 31464 38108 31476
rect 38063 31436 38108 31464
rect 38102 31424 38108 31436
rect 38160 31424 38166 31476
rect 38657 31467 38715 31473
rect 38657 31433 38669 31467
rect 38703 31464 38715 31467
rect 39850 31464 39856 31476
rect 38703 31436 39856 31464
rect 38703 31433 38715 31436
rect 38657 31427 38715 31433
rect 39850 31424 39856 31436
rect 39908 31424 39914 31476
rect 40310 31464 40316 31476
rect 40223 31436 40316 31464
rect 38838 31405 38844 31408
rect 38825 31399 38844 31405
rect 38825 31365 38837 31399
rect 38825 31359 38844 31365
rect 38838 31356 38844 31359
rect 38896 31356 38902 31408
rect 39022 31396 39028 31408
rect 38983 31368 39028 31396
rect 39022 31356 39028 31368
rect 39080 31356 39086 31408
rect 39482 31396 39488 31408
rect 39132 31368 39488 31396
rect 34992 31300 36400 31328
rect 33321 31291 33379 31297
rect 33597 31263 33655 31269
rect 33597 31229 33609 31263
rect 33643 31260 33655 31263
rect 33686 31260 33692 31272
rect 33643 31232 33692 31260
rect 33643 31229 33655 31232
rect 33597 31223 33655 31229
rect 33686 31220 33692 31232
rect 33744 31220 33750 31272
rect 35989 31263 36047 31269
rect 35989 31229 36001 31263
rect 36035 31229 36047 31263
rect 35989 31223 36047 31229
rect 33962 31084 33968 31136
rect 34020 31124 34026 31136
rect 35529 31127 35587 31133
rect 35529 31124 35541 31127
rect 34020 31096 35541 31124
rect 34020 31084 34026 31096
rect 35529 31093 35541 31096
rect 35575 31093 35587 31127
rect 35529 31087 35587 31093
rect 35802 31084 35808 31136
rect 35860 31124 35866 31136
rect 36004 31124 36032 31223
rect 36078 31220 36084 31272
rect 36136 31260 36142 31272
rect 36372 31260 36400 31300
rect 36446 31288 36452 31340
rect 36504 31328 36510 31340
rect 37461 31331 37519 31337
rect 37461 31328 37473 31331
rect 36504 31300 37473 31328
rect 36504 31288 36510 31300
rect 37461 31297 37473 31300
rect 37507 31328 37519 31331
rect 39132 31328 39160 31368
rect 39482 31356 39488 31368
rect 39540 31356 39546 31408
rect 40236 31405 40264 31436
rect 40310 31424 40316 31436
rect 40368 31464 40374 31476
rect 41322 31464 41328 31476
rect 40368 31436 41328 31464
rect 40368 31424 40374 31436
rect 41322 31424 41328 31436
rect 41380 31424 41386 31476
rect 45922 31424 45928 31476
rect 45980 31464 45986 31476
rect 46109 31467 46167 31473
rect 46109 31464 46121 31467
rect 45980 31436 46121 31464
rect 45980 31424 45986 31436
rect 46109 31433 46121 31436
rect 46155 31433 46167 31467
rect 48314 31464 48320 31476
rect 46109 31427 46167 31433
rect 46768 31436 48320 31464
rect 40221 31399 40279 31405
rect 40221 31365 40233 31399
rect 40267 31365 40279 31399
rect 40221 31359 40279 31365
rect 40451 31399 40509 31405
rect 40451 31365 40463 31399
rect 40497 31396 40509 31399
rect 40586 31396 40592 31408
rect 40497 31368 40592 31396
rect 40497 31365 40509 31368
rect 40451 31359 40509 31365
rect 40586 31356 40592 31368
rect 40644 31396 40650 31408
rect 41187 31399 41245 31405
rect 41187 31396 41199 31399
rect 40644 31368 41199 31396
rect 40644 31356 40650 31368
rect 41187 31365 41199 31368
rect 41233 31365 41245 31399
rect 41340 31396 41368 31424
rect 41417 31399 41475 31405
rect 41417 31396 41429 31399
rect 41340 31368 41429 31396
rect 41187 31359 41245 31365
rect 41417 31365 41429 31368
rect 41463 31365 41475 31399
rect 46014 31396 46020 31408
rect 45975 31368 46020 31396
rect 41417 31359 41475 31365
rect 46014 31356 46020 31368
rect 46072 31356 46078 31408
rect 37507 31300 39160 31328
rect 37507 31297 37519 31300
rect 37461 31291 37519 31297
rect 39298 31288 39304 31340
rect 39356 31328 39362 31340
rect 39758 31328 39764 31340
rect 39356 31300 39764 31328
rect 39356 31288 39362 31300
rect 39758 31288 39764 31300
rect 39816 31328 39822 31340
rect 40129 31331 40187 31337
rect 40129 31328 40141 31331
rect 39816 31300 40141 31328
rect 39816 31288 39822 31300
rect 40129 31297 40141 31300
rect 40175 31297 40187 31331
rect 40129 31291 40187 31297
rect 40313 31331 40371 31337
rect 40313 31297 40325 31331
rect 40359 31328 40371 31331
rect 40862 31328 40868 31340
rect 40359 31300 40868 31328
rect 40359 31297 40371 31300
rect 40313 31291 40371 31297
rect 39945 31263 40003 31269
rect 39945 31260 39957 31263
rect 36136 31232 36181 31260
rect 36372 31232 39957 31260
rect 36136 31220 36142 31232
rect 39945 31229 39957 31232
rect 39991 31229 40003 31263
rect 39945 31223 40003 31229
rect 40034 31220 40040 31272
rect 40092 31260 40098 31272
rect 40328 31260 40356 31291
rect 40862 31288 40868 31300
rect 40920 31328 40926 31340
rect 41325 31331 41383 31337
rect 41325 31328 41337 31331
rect 40920 31300 41337 31328
rect 40920 31288 40926 31300
rect 41325 31297 41337 31300
rect 41371 31297 41383 31331
rect 41506 31328 41512 31340
rect 41467 31300 41512 31328
rect 41325 31291 41383 31297
rect 41506 31288 41512 31300
rect 41564 31288 41570 31340
rect 43346 31328 43352 31340
rect 43307 31300 43352 31328
rect 43346 31288 43352 31300
rect 43404 31328 43410 31340
rect 43714 31328 43720 31340
rect 43404 31300 43720 31328
rect 43404 31288 43410 31300
rect 43714 31288 43720 31300
rect 43772 31288 43778 31340
rect 44082 31328 44088 31340
rect 44043 31300 44088 31328
rect 44082 31288 44088 31300
rect 44140 31288 44146 31340
rect 45186 31328 45192 31340
rect 45147 31300 45192 31328
rect 45186 31288 45192 31300
rect 45244 31328 45250 31340
rect 46768 31328 46796 31436
rect 48314 31424 48320 31436
rect 48372 31424 48378 31476
rect 50709 31467 50767 31473
rect 50709 31433 50721 31467
rect 50755 31433 50767 31467
rect 50709 31427 50767 31433
rect 50893 31467 50951 31473
rect 50893 31433 50905 31467
rect 50939 31464 50951 31467
rect 50982 31464 50988 31476
rect 50939 31436 50988 31464
rect 50939 31433 50951 31436
rect 50893 31427 50951 31433
rect 46842 31356 46848 31408
rect 46900 31396 46906 31408
rect 47670 31396 47676 31408
rect 46900 31368 47676 31396
rect 46900 31356 46906 31368
rect 47670 31356 47676 31368
rect 47728 31356 47734 31408
rect 48332 31396 48360 31424
rect 50724 31396 50752 31427
rect 50982 31424 50988 31436
rect 51040 31424 51046 31476
rect 51721 31467 51779 31473
rect 51721 31433 51733 31467
rect 51767 31464 51779 31467
rect 52638 31464 52644 31476
rect 51767 31436 52644 31464
rect 51767 31433 51779 31436
rect 51721 31427 51779 31433
rect 52638 31424 52644 31436
rect 52696 31464 52702 31476
rect 55217 31467 55275 31473
rect 55217 31464 55229 31467
rect 52696 31436 55229 31464
rect 52696 31424 52702 31436
rect 55217 31433 55229 31436
rect 55263 31433 55275 31467
rect 55217 31427 55275 31433
rect 56413 31467 56471 31473
rect 56413 31433 56425 31467
rect 56459 31433 56471 31467
rect 56413 31427 56471 31433
rect 51902 31396 51908 31408
rect 48332 31368 49188 31396
rect 50724 31368 51028 31396
rect 46934 31328 46940 31340
rect 45244 31300 46796 31328
rect 46895 31300 46940 31328
rect 45244 31288 45250 31300
rect 46934 31288 46940 31300
rect 46992 31288 46998 31340
rect 47121 31331 47179 31337
rect 47121 31297 47133 31331
rect 47167 31297 47179 31331
rect 47121 31291 47179 31297
rect 40092 31232 40356 31260
rect 40589 31263 40647 31269
rect 40092 31220 40098 31232
rect 40589 31229 40601 31263
rect 40635 31229 40647 31263
rect 40589 31223 40647 31229
rect 41049 31263 41107 31269
rect 41049 31229 41061 31263
rect 41095 31260 41107 31263
rect 42886 31260 42892 31272
rect 41095 31232 42892 31260
rect 41095 31229 41107 31232
rect 41049 31223 41107 31229
rect 36096 31192 36124 31220
rect 36998 31192 37004 31204
rect 36096 31164 37004 31192
rect 36998 31152 37004 31164
rect 37056 31152 37062 31204
rect 39022 31192 39028 31204
rect 37384 31164 39028 31192
rect 36725 31127 36783 31133
rect 36725 31124 36737 31127
rect 35860 31096 36737 31124
rect 35860 31084 35866 31096
rect 36725 31093 36737 31096
rect 36771 31124 36783 31127
rect 37384 31124 37412 31164
rect 39022 31152 39028 31164
rect 39080 31152 39086 31204
rect 40604 31192 40632 31223
rect 42886 31220 42892 31232
rect 42944 31220 42950 31272
rect 42978 31220 42984 31272
rect 43036 31260 43042 31272
rect 44634 31260 44640 31272
rect 43036 31232 44640 31260
rect 43036 31220 43042 31232
rect 44634 31220 44640 31232
rect 44692 31260 44698 31272
rect 44913 31263 44971 31269
rect 44913 31260 44925 31263
rect 44692 31232 44925 31260
rect 44692 31220 44698 31232
rect 44913 31229 44925 31232
rect 44959 31229 44971 31263
rect 44913 31223 44971 31229
rect 45925 31263 45983 31269
rect 45925 31229 45937 31263
rect 45971 31260 45983 31263
rect 46198 31260 46204 31272
rect 45971 31232 46204 31260
rect 45971 31229 45983 31232
rect 45925 31223 45983 31229
rect 46198 31220 46204 31232
rect 46256 31260 46262 31272
rect 47136 31260 47164 31291
rect 46256 31232 47164 31260
rect 47688 31260 47716 31356
rect 47765 31331 47823 31337
rect 47765 31297 47777 31331
rect 47811 31328 47823 31331
rect 48314 31328 48320 31340
rect 47811 31300 48320 31328
rect 47811 31297 47823 31300
rect 47765 31291 47823 31297
rect 48314 31288 48320 31300
rect 48372 31288 48378 31340
rect 49160 31337 49188 31368
rect 50798 31337 50804 31340
rect 49145 31331 49203 31337
rect 49145 31297 49157 31331
rect 49191 31297 49203 31331
rect 49145 31291 49203 31297
rect 49329 31331 49387 31337
rect 49329 31297 49341 31331
rect 49375 31328 49387 31331
rect 50768 31331 50804 31337
rect 49375 31300 50384 31328
rect 49375 31297 49387 31300
rect 49329 31291 49387 31297
rect 47857 31263 47915 31269
rect 47857 31260 47869 31263
rect 47688 31232 47869 31260
rect 46256 31220 46262 31232
rect 47857 31229 47869 31232
rect 47903 31229 47915 31263
rect 48958 31260 48964 31272
rect 48919 31232 48964 31260
rect 47857 31223 47915 31229
rect 42426 31192 42432 31204
rect 40604 31164 42432 31192
rect 42426 31152 42432 31164
rect 42484 31152 42490 31204
rect 42702 31192 42708 31204
rect 42663 31164 42708 31192
rect 42702 31152 42708 31164
rect 42760 31152 42766 31204
rect 43162 31192 43168 31204
rect 43123 31164 43168 31192
rect 43162 31152 43168 31164
rect 43220 31152 43226 31204
rect 46477 31195 46535 31201
rect 46477 31161 46489 31195
rect 46523 31192 46535 31195
rect 47210 31192 47216 31204
rect 46523 31164 47216 31192
rect 46523 31161 46535 31164
rect 46477 31155 46535 31161
rect 47210 31152 47216 31164
rect 47268 31152 47274 31204
rect 36771 31096 37412 31124
rect 36771 31093 36783 31096
rect 36725 31087 36783 31093
rect 37458 31084 37464 31136
rect 37516 31124 37522 31136
rect 37553 31127 37611 31133
rect 37553 31124 37565 31127
rect 37516 31096 37565 31124
rect 37516 31084 37522 31096
rect 37553 31093 37565 31096
rect 37599 31093 37611 31127
rect 37553 31087 37611 31093
rect 38746 31084 38752 31136
rect 38804 31124 38810 31136
rect 38841 31127 38899 31133
rect 38841 31124 38853 31127
rect 38804 31096 38853 31124
rect 38804 31084 38810 31096
rect 38841 31093 38853 31096
rect 38887 31093 38899 31127
rect 38841 31087 38899 31093
rect 41693 31127 41751 31133
rect 41693 31093 41705 31127
rect 41739 31124 41751 31127
rect 41782 31124 41788 31136
rect 41739 31096 41788 31124
rect 41739 31093 41751 31096
rect 41693 31087 41751 31093
rect 41782 31084 41788 31096
rect 41840 31084 41846 31136
rect 43438 31084 43444 31136
rect 43496 31124 43502 31136
rect 43993 31127 44051 31133
rect 43993 31124 44005 31127
rect 43496 31096 44005 31124
rect 43496 31084 43502 31096
rect 43993 31093 44005 31096
rect 44039 31093 44051 31127
rect 46934 31124 46940 31136
rect 46895 31096 46940 31124
rect 43993 31087 44051 31093
rect 46934 31084 46940 31096
rect 46992 31084 46998 31136
rect 47026 31084 47032 31136
rect 47084 31124 47090 31136
rect 47765 31127 47823 31133
rect 47765 31124 47777 31127
rect 47084 31096 47777 31124
rect 47084 31084 47090 31096
rect 47765 31093 47777 31096
rect 47811 31093 47823 31127
rect 47872 31124 47900 31223
rect 48958 31220 48964 31232
rect 49016 31220 49022 31272
rect 50249 31263 50307 31269
rect 50249 31229 50261 31263
rect 50295 31229 50307 31263
rect 50249 31223 50307 31229
rect 48133 31195 48191 31201
rect 48133 31161 48145 31195
rect 48179 31192 48191 31195
rect 48406 31192 48412 31204
rect 48179 31164 48412 31192
rect 48179 31161 48191 31164
rect 48133 31155 48191 31161
rect 48406 31152 48412 31164
rect 48464 31192 48470 31204
rect 50264 31192 50292 31223
rect 50356 31204 50384 31300
rect 50768 31297 50780 31331
rect 50768 31291 50804 31297
rect 50798 31288 50804 31291
rect 50856 31288 50862 31340
rect 51000 31328 51028 31368
rect 51368 31368 51908 31396
rect 51368 31328 51396 31368
rect 51902 31356 51908 31368
rect 51960 31356 51966 31408
rect 53558 31396 53564 31408
rect 53116 31368 53564 31396
rect 51534 31328 51540 31340
rect 51000 31300 51396 31328
rect 51495 31300 51540 31328
rect 51534 31288 51540 31300
rect 51592 31288 51598 31340
rect 51813 31331 51871 31337
rect 51813 31297 51825 31331
rect 51859 31328 51871 31331
rect 53116 31328 53144 31368
rect 53558 31356 53564 31368
rect 53616 31356 53622 31408
rect 54110 31356 54116 31408
rect 54168 31396 54174 31408
rect 54205 31399 54263 31405
rect 54205 31396 54217 31399
rect 54168 31368 54217 31396
rect 54168 31356 54174 31368
rect 54205 31365 54217 31368
rect 54251 31396 54263 31399
rect 55861 31399 55919 31405
rect 54251 31368 55812 31396
rect 54251 31365 54263 31368
rect 54205 31359 54263 31365
rect 51859 31300 53144 31328
rect 53193 31331 53251 31337
rect 51859 31297 51871 31300
rect 51813 31291 51871 31297
rect 53193 31297 53205 31331
rect 53239 31328 53251 31331
rect 53742 31328 53748 31340
rect 53239 31300 53748 31328
rect 53239 31297 53251 31300
rect 53193 31291 53251 31297
rect 53742 31288 53748 31300
rect 53800 31328 53806 31340
rect 54294 31328 54300 31340
rect 53800 31300 54300 31328
rect 53800 31288 53806 31300
rect 54294 31288 54300 31300
rect 54352 31288 54358 31340
rect 54478 31328 54484 31340
rect 54439 31300 54484 31328
rect 54478 31288 54484 31300
rect 54536 31288 54542 31340
rect 54570 31288 54576 31340
rect 54628 31328 54634 31340
rect 55030 31328 55036 31340
rect 54628 31300 55036 31328
rect 54628 31288 54634 31300
rect 55030 31288 55036 31300
rect 55088 31288 55094 31340
rect 55784 31328 55812 31368
rect 55861 31365 55873 31399
rect 55907 31396 55919 31399
rect 56318 31396 56324 31408
rect 55907 31368 56324 31396
rect 55907 31365 55919 31368
rect 55861 31359 55919 31365
rect 56318 31356 56324 31368
rect 56376 31356 56382 31408
rect 56134 31328 56140 31340
rect 55784 31300 55996 31328
rect 56095 31300 56140 31328
rect 52273 31263 52331 31269
rect 52273 31260 52285 31263
rect 51046 31232 52285 31260
rect 48464 31164 50292 31192
rect 48464 31152 48470 31164
rect 50338 31152 50344 31204
rect 50396 31192 50402 31204
rect 50396 31164 50441 31192
rect 50396 31152 50402 31164
rect 49602 31124 49608 31136
rect 47872 31096 49608 31124
rect 47765 31087 47823 31093
rect 49602 31084 49608 31096
rect 49660 31084 49666 31136
rect 49878 31084 49884 31136
rect 49936 31124 49942 31136
rect 51046 31124 51074 31232
rect 52273 31229 52285 31232
rect 52319 31229 52331 31263
rect 54110 31260 54116 31272
rect 54071 31232 54116 31260
rect 52273 31223 52331 31229
rect 54110 31220 54116 31232
rect 54168 31260 54174 31272
rect 54386 31260 54392 31272
rect 54168 31232 54392 31260
rect 54168 31220 54174 31232
rect 54386 31220 54392 31232
rect 54444 31220 54450 31272
rect 55582 31220 55588 31272
rect 55640 31260 55646 31272
rect 55769 31263 55827 31269
rect 55769 31260 55781 31263
rect 55640 31232 55781 31260
rect 55640 31220 55646 31232
rect 55769 31229 55781 31232
rect 55815 31229 55827 31263
rect 55968 31260 55996 31300
rect 56134 31288 56140 31300
rect 56192 31288 56198 31340
rect 56428 31328 56456 31427
rect 56778 31356 56784 31408
rect 56836 31396 56842 31408
rect 56836 31368 57008 31396
rect 56836 31356 56842 31368
rect 56980 31337 57008 31368
rect 57054 31356 57060 31408
rect 57112 31396 57118 31408
rect 57112 31368 57284 31396
rect 57112 31356 57118 31368
rect 57256 31337 57284 31368
rect 56873 31331 56931 31337
rect 56873 31328 56885 31331
rect 56428 31300 56885 31328
rect 56873 31297 56885 31300
rect 56919 31297 56931 31331
rect 56873 31291 56931 31297
rect 56965 31331 57023 31337
rect 56965 31297 56977 31331
rect 57011 31297 57023 31331
rect 56965 31291 57023 31297
rect 57149 31331 57207 31337
rect 57149 31297 57161 31331
rect 57195 31297 57207 31331
rect 57149 31291 57207 31297
rect 57241 31331 57299 31337
rect 57241 31297 57253 31331
rect 57287 31297 57299 31331
rect 57241 31291 57299 31297
rect 58345 31331 58403 31337
rect 58345 31297 58357 31331
rect 58391 31328 58403 31331
rect 58526 31328 58532 31340
rect 58391 31300 58532 31328
rect 58391 31297 58403 31300
rect 58345 31291 58403 31297
rect 56229 31263 56287 31269
rect 56229 31260 56241 31263
rect 55968 31232 56241 31260
rect 55769 31223 55827 31229
rect 56229 31229 56241 31232
rect 56275 31260 56287 31263
rect 57164 31260 57192 31291
rect 58526 31288 58532 31300
rect 58584 31288 58590 31340
rect 57882 31260 57888 31272
rect 56275 31232 57888 31260
rect 56275 31229 56287 31232
rect 56229 31223 56287 31229
rect 57882 31220 57888 31232
rect 57940 31220 57946 31272
rect 58066 31260 58072 31272
rect 58027 31232 58072 31260
rect 58066 31220 58072 31232
rect 58124 31220 58130 31272
rect 57606 31152 57612 31204
rect 57664 31192 57670 31204
rect 58253 31195 58311 31201
rect 58253 31192 58265 31195
rect 57664 31164 58265 31192
rect 57664 31152 57670 31164
rect 58253 31161 58265 31164
rect 58299 31161 58311 31195
rect 58253 31155 58311 31161
rect 51350 31124 51356 31136
rect 49936 31096 51074 31124
rect 51311 31096 51356 31124
rect 49936 31084 49942 31096
rect 51350 31084 51356 31096
rect 51408 31084 51414 31136
rect 52270 31084 52276 31136
rect 52328 31124 52334 31136
rect 53009 31127 53067 31133
rect 53009 31124 53021 31127
rect 52328 31096 53021 31124
rect 52328 31084 52334 31096
rect 53009 31093 53021 31096
rect 53055 31124 53067 31127
rect 53374 31124 53380 31136
rect 53055 31096 53380 31124
rect 53055 31093 53067 31096
rect 53009 31087 53067 31093
rect 53374 31084 53380 31096
rect 53432 31084 53438 31136
rect 54754 31124 54760 31136
rect 54715 31096 54760 31124
rect 54754 31084 54760 31096
rect 54812 31084 54818 31136
rect 57146 31084 57152 31136
rect 57204 31124 57210 31136
rect 57425 31127 57483 31133
rect 57425 31124 57437 31127
rect 57204 31096 57437 31124
rect 57204 31084 57210 31096
rect 57425 31093 57437 31096
rect 57471 31093 57483 31127
rect 57425 31087 57483 31093
rect 57790 31084 57796 31136
rect 57848 31124 57854 31136
rect 58161 31127 58219 31133
rect 58161 31124 58173 31127
rect 57848 31096 58173 31124
rect 57848 31084 57854 31096
rect 58161 31093 58173 31096
rect 58207 31093 58219 31127
rect 58161 31087 58219 31093
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 33686 30920 33692 30932
rect 33647 30892 33692 30920
rect 33686 30880 33692 30892
rect 33744 30880 33750 30932
rect 38746 30880 38752 30932
rect 38804 30920 38810 30932
rect 39117 30923 39175 30929
rect 39117 30920 39129 30923
rect 38804 30892 39129 30920
rect 38804 30880 38810 30892
rect 39117 30889 39129 30892
rect 39163 30889 39175 30923
rect 39117 30883 39175 30889
rect 39301 30923 39359 30929
rect 39301 30889 39313 30923
rect 39347 30920 39359 30923
rect 40402 30920 40408 30932
rect 39347 30892 40408 30920
rect 39347 30889 39359 30892
rect 39301 30883 39359 30889
rect 40402 30880 40408 30892
rect 40460 30880 40466 30932
rect 43257 30923 43315 30929
rect 43257 30889 43269 30923
rect 43303 30920 43315 30923
rect 44266 30920 44272 30932
rect 43303 30892 44272 30920
rect 43303 30889 43315 30892
rect 43257 30883 43315 30889
rect 44266 30880 44272 30892
rect 44324 30880 44330 30932
rect 46566 30880 46572 30932
rect 46624 30920 46630 30932
rect 49421 30923 49479 30929
rect 46624 30892 48912 30920
rect 46624 30880 46630 30892
rect 33870 30812 33876 30864
rect 33928 30852 33934 30864
rect 38197 30855 38255 30861
rect 33928 30824 35940 30852
rect 33928 30812 33934 30824
rect 29454 30744 29460 30796
rect 29512 30784 29518 30796
rect 29825 30787 29883 30793
rect 29825 30784 29837 30787
rect 29512 30756 29837 30784
rect 29512 30744 29518 30756
rect 29825 30753 29837 30756
rect 29871 30753 29883 30787
rect 29825 30747 29883 30753
rect 34790 30744 34796 30796
rect 34848 30784 34854 30796
rect 35342 30784 35348 30796
rect 34848 30756 35348 30784
rect 34848 30744 34854 30756
rect 35342 30744 35348 30756
rect 35400 30784 35406 30796
rect 35437 30787 35495 30793
rect 35437 30784 35449 30787
rect 35400 30756 35449 30784
rect 35400 30744 35406 30756
rect 35437 30753 35449 30756
rect 35483 30753 35495 30787
rect 35912 30784 35940 30824
rect 38197 30821 38209 30855
rect 38243 30852 38255 30855
rect 39390 30852 39396 30864
rect 38243 30824 39396 30852
rect 38243 30821 38255 30824
rect 38197 30815 38255 30821
rect 39390 30812 39396 30824
rect 39448 30812 39454 30864
rect 45925 30855 45983 30861
rect 45925 30821 45937 30855
rect 45971 30852 45983 30855
rect 48884 30852 48912 30892
rect 49421 30889 49433 30923
rect 49467 30920 49479 30923
rect 51534 30920 51540 30932
rect 49467 30892 51540 30920
rect 49467 30889 49479 30892
rect 49421 30883 49479 30889
rect 51534 30880 51540 30892
rect 51592 30880 51598 30932
rect 53469 30923 53527 30929
rect 53469 30889 53481 30923
rect 53515 30920 53527 30923
rect 55858 30920 55864 30932
rect 53515 30892 55864 30920
rect 53515 30889 53527 30892
rect 53469 30883 53527 30889
rect 50982 30852 50988 30864
rect 45971 30824 48820 30852
rect 48884 30824 50988 30852
rect 45971 30821 45983 30824
rect 45925 30815 45983 30821
rect 40037 30787 40095 30793
rect 40037 30784 40049 30787
rect 35912 30756 40049 30784
rect 35437 30747 35495 30753
rect 40037 30753 40049 30756
rect 40083 30753 40095 30787
rect 40037 30747 40095 30753
rect 41509 30787 41567 30793
rect 41509 30753 41521 30787
rect 41555 30784 41567 30787
rect 43346 30784 43352 30796
rect 41555 30756 43352 30784
rect 41555 30753 41567 30756
rect 41509 30747 41567 30753
rect 43346 30744 43352 30756
rect 43404 30744 43410 30796
rect 47397 30787 47455 30793
rect 47397 30784 47409 30787
rect 46492 30756 47409 30784
rect 1857 30719 1915 30725
rect 1857 30685 1869 30719
rect 1903 30716 1915 30719
rect 1903 30688 2452 30716
rect 1903 30685 1915 30688
rect 1857 30679 1915 30685
rect 2424 30592 2452 30688
rect 31846 30676 31852 30728
rect 31904 30716 31910 30728
rect 33045 30719 33103 30725
rect 31904 30688 31949 30716
rect 31904 30676 31910 30688
rect 33045 30685 33057 30719
rect 33091 30685 33103 30719
rect 33045 30679 33103 30685
rect 33873 30719 33931 30725
rect 33873 30685 33885 30719
rect 33919 30716 33931 30719
rect 33962 30716 33968 30728
rect 33919 30688 33968 30716
rect 33919 30685 33931 30688
rect 33873 30679 33931 30685
rect 30834 30608 30840 30660
rect 30892 30608 30898 30660
rect 31573 30651 31631 30657
rect 31573 30617 31585 30651
rect 31619 30648 31631 30651
rect 31662 30648 31668 30660
rect 31619 30620 31668 30648
rect 31619 30617 31631 30620
rect 31573 30611 31631 30617
rect 31662 30608 31668 30620
rect 31720 30608 31726 30660
rect 33060 30648 33088 30679
rect 33962 30676 33968 30688
rect 34020 30676 34026 30728
rect 34146 30676 34152 30728
rect 34204 30716 34210 30728
rect 36449 30719 36507 30725
rect 36449 30716 36461 30719
rect 34204 30688 36461 30716
rect 34204 30676 34210 30688
rect 36449 30685 36461 30688
rect 36495 30685 36507 30719
rect 36449 30679 36507 30685
rect 39758 30676 39764 30728
rect 39816 30716 39822 30728
rect 40221 30719 40279 30725
rect 40221 30716 40233 30719
rect 39816 30688 40233 30716
rect 39816 30676 39822 30688
rect 40221 30685 40233 30688
rect 40267 30685 40279 30719
rect 40402 30716 40408 30728
rect 40363 30688 40408 30716
rect 40221 30679 40279 30685
rect 40402 30676 40408 30688
rect 40460 30676 40466 30728
rect 40681 30719 40739 30725
rect 40681 30685 40693 30719
rect 40727 30716 40739 30719
rect 40770 30716 40776 30728
rect 40727 30688 40776 30716
rect 40727 30685 40739 30688
rect 40681 30679 40739 30685
rect 40770 30676 40776 30688
rect 40828 30716 40834 30728
rect 41322 30716 41328 30728
rect 40828 30688 41328 30716
rect 40828 30676 40834 30688
rect 41322 30676 41328 30688
rect 41380 30676 41386 30728
rect 43070 30676 43076 30728
rect 43128 30716 43134 30728
rect 43809 30719 43867 30725
rect 43809 30716 43821 30719
rect 43128 30688 43821 30716
rect 43128 30676 43134 30688
rect 43809 30685 43821 30688
rect 43855 30685 43867 30719
rect 43809 30679 43867 30685
rect 43898 30676 43904 30728
rect 43956 30716 43962 30728
rect 43993 30719 44051 30725
rect 43993 30716 44005 30719
rect 43956 30688 44005 30716
rect 43956 30676 43962 30688
rect 43993 30685 44005 30688
rect 44039 30685 44051 30719
rect 43993 30679 44051 30685
rect 45465 30719 45523 30725
rect 45465 30685 45477 30719
rect 45511 30685 45523 30719
rect 45465 30679 45523 30685
rect 45741 30719 45799 30725
rect 45741 30685 45753 30719
rect 45787 30716 45799 30719
rect 45922 30716 45928 30728
rect 45787 30688 45928 30716
rect 45787 30685 45799 30688
rect 45741 30679 45799 30685
rect 35253 30651 35311 30657
rect 33060 30620 34928 30648
rect 1670 30580 1676 30592
rect 1631 30552 1676 30580
rect 1670 30540 1676 30552
rect 1728 30540 1734 30592
rect 2406 30580 2412 30592
rect 2367 30552 2412 30580
rect 2406 30540 2412 30552
rect 2464 30540 2470 30592
rect 33229 30583 33287 30589
rect 33229 30549 33241 30583
rect 33275 30580 33287 30583
rect 34790 30580 34796 30592
rect 33275 30552 34796 30580
rect 33275 30549 33287 30552
rect 33229 30543 33287 30549
rect 34790 30540 34796 30552
rect 34848 30540 34854 30592
rect 34900 30589 34928 30620
rect 35253 30617 35265 30651
rect 35299 30648 35311 30651
rect 36170 30648 36176 30660
rect 35299 30620 36176 30648
rect 35299 30617 35311 30620
rect 35253 30611 35311 30617
rect 36170 30608 36176 30620
rect 36228 30648 36234 30660
rect 36354 30648 36360 30660
rect 36228 30620 36360 30648
rect 36228 30608 36234 30620
rect 36354 30608 36360 30620
rect 36412 30608 36418 30660
rect 36725 30651 36783 30657
rect 36725 30617 36737 30651
rect 36771 30617 36783 30651
rect 36725 30611 36783 30617
rect 34885 30583 34943 30589
rect 34885 30549 34897 30583
rect 34931 30549 34943 30583
rect 34885 30543 34943 30549
rect 35158 30540 35164 30592
rect 35216 30580 35222 30592
rect 35345 30583 35403 30589
rect 35345 30580 35357 30583
rect 35216 30552 35357 30580
rect 35216 30540 35222 30552
rect 35345 30549 35357 30552
rect 35391 30580 35403 30583
rect 35802 30580 35808 30592
rect 35391 30552 35808 30580
rect 35391 30549 35403 30552
rect 35345 30543 35403 30549
rect 35802 30540 35808 30552
rect 35860 30540 35866 30592
rect 36446 30540 36452 30592
rect 36504 30580 36510 30592
rect 36740 30580 36768 30611
rect 37458 30608 37464 30660
rect 37516 30608 37522 30660
rect 38930 30648 38936 30660
rect 38891 30620 38936 30648
rect 38930 30608 38936 30620
rect 38988 30608 38994 30660
rect 40034 30608 40040 30660
rect 40092 30648 40098 30660
rect 40310 30648 40316 30660
rect 40092 30620 40316 30648
rect 40092 30608 40098 30620
rect 40310 30608 40316 30620
rect 40368 30608 40374 30660
rect 40494 30608 40500 30660
rect 40552 30657 40558 30660
rect 40552 30651 40581 30657
rect 40569 30617 40581 30651
rect 41782 30648 41788 30660
rect 41743 30620 41788 30648
rect 40552 30611 40581 30617
rect 40552 30608 40558 30611
rect 41782 30608 41788 30620
rect 41840 30608 41846 30660
rect 43438 30648 43444 30660
rect 43010 30620 43444 30648
rect 43438 30608 43444 30620
rect 43496 30608 43502 30660
rect 43714 30608 43720 30660
rect 43772 30648 43778 30660
rect 45278 30648 45284 30660
rect 43772 30620 45284 30648
rect 43772 30608 43778 30620
rect 45278 30608 45284 30620
rect 45336 30648 45342 30660
rect 45480 30648 45508 30679
rect 45922 30676 45928 30688
rect 45980 30676 45986 30728
rect 46106 30676 46112 30728
rect 46164 30716 46170 30728
rect 46492 30725 46520 30756
rect 47397 30753 47409 30756
rect 47443 30753 47455 30787
rect 48406 30784 48412 30796
rect 47397 30747 47455 30753
rect 47780 30756 48412 30784
rect 46385 30719 46443 30725
rect 46385 30716 46397 30719
rect 46164 30688 46397 30716
rect 46164 30676 46170 30688
rect 46385 30685 46397 30688
rect 46431 30685 46443 30719
rect 46385 30679 46443 30685
rect 46477 30719 46535 30725
rect 46477 30685 46489 30719
rect 46523 30685 46535 30719
rect 46477 30679 46535 30685
rect 46566 30676 46572 30728
rect 46624 30716 46630 30728
rect 46661 30719 46719 30725
rect 46661 30716 46673 30719
rect 46624 30688 46673 30716
rect 46624 30676 46630 30688
rect 46661 30685 46673 30688
rect 46707 30685 46719 30719
rect 46661 30679 46719 30685
rect 46750 30676 46756 30728
rect 46808 30716 46814 30728
rect 47578 30716 47584 30728
rect 46808 30688 46853 30716
rect 47539 30688 47584 30716
rect 46808 30676 46814 30688
rect 47578 30676 47584 30688
rect 47636 30676 47642 30728
rect 47673 30719 47731 30725
rect 47673 30685 47685 30719
rect 47719 30716 47731 30719
rect 47780 30716 47808 30756
rect 48406 30744 48412 30756
rect 48464 30744 48470 30796
rect 48792 30793 48820 30824
rect 50982 30812 50988 30824
rect 51040 30852 51046 30864
rect 53484 30852 53512 30883
rect 55858 30880 55864 30892
rect 55916 30880 55922 30932
rect 57517 30923 57575 30929
rect 57517 30889 57529 30923
rect 57563 30920 57575 30923
rect 57606 30920 57612 30932
rect 57563 30892 57612 30920
rect 57563 30889 57575 30892
rect 57517 30883 57575 30889
rect 57606 30880 57612 30892
rect 57664 30880 57670 30932
rect 51040 30824 53512 30852
rect 51040 30812 51046 30824
rect 54018 30812 54024 30864
rect 54076 30852 54082 30864
rect 54076 30824 54156 30852
rect 54076 30812 54082 30824
rect 48777 30787 48835 30793
rect 48777 30753 48789 30787
rect 48823 30753 48835 30787
rect 48777 30747 48835 30753
rect 48961 30787 49019 30793
rect 48961 30753 48973 30787
rect 49007 30784 49019 30787
rect 50338 30784 50344 30796
rect 49007 30756 50344 30784
rect 49007 30753 49019 30756
rect 48961 30747 49019 30753
rect 50338 30744 50344 30756
rect 50396 30784 50402 30796
rect 50798 30784 50804 30796
rect 50396 30756 50804 30784
rect 50396 30744 50402 30756
rect 50798 30744 50804 30756
rect 50856 30784 50862 30796
rect 51442 30784 51448 30796
rect 50856 30756 51448 30784
rect 50856 30744 50862 30756
rect 47719 30688 47808 30716
rect 47719 30685 47731 30688
rect 47673 30679 47731 30685
rect 47854 30676 47860 30728
rect 47912 30725 47918 30728
rect 47912 30719 47941 30725
rect 47929 30685 47941 30719
rect 48038 30716 48044 30728
rect 47999 30688 48044 30716
rect 47912 30679 47941 30685
rect 47912 30676 47918 30679
rect 48038 30676 48044 30688
rect 48096 30676 48102 30728
rect 49050 30716 49056 30728
rect 49011 30688 49056 30716
rect 49050 30676 49056 30688
rect 49108 30676 49114 30728
rect 51000 30725 51028 30756
rect 51442 30744 51448 30756
rect 51500 30744 51506 30796
rect 52454 30784 52460 30796
rect 52415 30756 52460 30784
rect 52454 30744 52460 30756
rect 52512 30784 52518 30796
rect 52730 30784 52736 30796
rect 52512 30756 52736 30784
rect 52512 30744 52518 30756
rect 52730 30744 52736 30756
rect 52788 30744 52794 30796
rect 54128 30784 54156 30824
rect 54294 30812 54300 30864
rect 54352 30812 54358 30864
rect 54570 30812 54576 30864
rect 54628 30852 54634 30864
rect 54628 30824 55812 30852
rect 54628 30812 54634 30824
rect 54205 30787 54263 30793
rect 54205 30784 54217 30787
rect 54128 30756 54217 30784
rect 54205 30753 54217 30756
rect 54251 30753 54263 30787
rect 54312 30784 54340 30812
rect 54312 30756 55628 30784
rect 54205 30747 54263 30753
rect 50709 30719 50767 30725
rect 50709 30685 50721 30719
rect 50755 30685 50767 30719
rect 50709 30679 50767 30685
rect 50985 30719 51043 30725
rect 50985 30685 50997 30719
rect 51031 30685 51043 30719
rect 51166 30716 51172 30728
rect 51127 30688 51172 30716
rect 50985 30679 51043 30685
rect 45336 30620 45508 30648
rect 47765 30651 47823 30657
rect 45336 30608 45342 30620
rect 47765 30617 47777 30651
rect 47811 30617 47823 30651
rect 47765 30611 47823 30617
rect 36504 30552 36768 30580
rect 36504 30540 36510 30552
rect 38838 30540 38844 30592
rect 38896 30580 38902 30592
rect 39133 30583 39191 30589
rect 39133 30580 39145 30583
rect 38896 30552 39145 30580
rect 38896 30540 38902 30552
rect 39133 30549 39145 30552
rect 39179 30549 39191 30583
rect 44174 30580 44180 30592
rect 44135 30552 44180 30580
rect 39133 30543 39191 30549
rect 44174 30540 44180 30552
rect 44232 30540 44238 30592
rect 45557 30583 45615 30589
rect 45557 30549 45569 30583
rect 45603 30580 45615 30583
rect 46014 30580 46020 30592
rect 45603 30552 46020 30580
rect 45603 30549 45615 30552
rect 45557 30543 45615 30549
rect 46014 30540 46020 30552
rect 46072 30580 46078 30592
rect 46842 30580 46848 30592
rect 46072 30552 46848 30580
rect 46072 30540 46078 30552
rect 46842 30540 46848 30552
rect 46900 30540 46906 30592
rect 46937 30583 46995 30589
rect 46937 30549 46949 30583
rect 46983 30580 46995 30583
rect 47578 30580 47584 30592
rect 46983 30552 47584 30580
rect 46983 30549 46995 30552
rect 46937 30543 46995 30549
rect 47578 30540 47584 30552
rect 47636 30540 47642 30592
rect 47670 30540 47676 30592
rect 47728 30580 47734 30592
rect 47781 30580 47809 30611
rect 48130 30608 48136 30660
rect 48188 30648 48194 30660
rect 49694 30648 49700 30660
rect 48188 30620 49700 30648
rect 48188 30608 48194 30620
rect 49694 30608 49700 30620
rect 49752 30608 49758 30660
rect 50614 30608 50620 30660
rect 50672 30648 50678 30660
rect 50724 30648 50752 30679
rect 51166 30676 51172 30688
rect 51224 30676 51230 30728
rect 51626 30716 51632 30728
rect 51276 30688 51632 30716
rect 51276 30648 51304 30688
rect 51626 30676 51632 30688
rect 51684 30676 51690 30728
rect 52546 30716 52552 30728
rect 52507 30688 52552 30716
rect 52546 30676 52552 30688
rect 52604 30716 52610 30728
rect 54297 30719 54355 30725
rect 54297 30716 54309 30719
rect 52604 30688 54309 30716
rect 52604 30676 52610 30688
rect 54297 30685 54309 30688
rect 54343 30716 54355 30719
rect 54478 30716 54484 30728
rect 54343 30688 54484 30716
rect 54343 30685 54355 30688
rect 54297 30679 54355 30685
rect 54478 30676 54484 30688
rect 54536 30676 54542 30728
rect 54754 30676 54760 30728
rect 54812 30716 54818 30728
rect 55600 30725 55628 30756
rect 55784 30725 55812 30824
rect 57241 30787 57299 30793
rect 57241 30753 57253 30787
rect 57287 30784 57299 30787
rect 57330 30784 57336 30796
rect 57287 30756 57336 30784
rect 57287 30753 57299 30756
rect 57241 30747 57299 30753
rect 57330 30744 57336 30756
rect 57388 30784 57394 30796
rect 58434 30784 58440 30796
rect 57388 30756 58440 30784
rect 57388 30744 57394 30756
rect 58434 30744 58440 30756
rect 58492 30744 58498 30796
rect 55493 30719 55551 30725
rect 55493 30716 55505 30719
rect 54812 30688 55505 30716
rect 54812 30676 54818 30688
rect 55493 30685 55505 30688
rect 55539 30685 55551 30719
rect 55493 30679 55551 30685
rect 55585 30719 55643 30725
rect 55585 30685 55597 30719
rect 55631 30685 55643 30719
rect 55585 30679 55643 30685
rect 55769 30719 55827 30725
rect 55769 30685 55781 30719
rect 55815 30685 55827 30719
rect 55769 30679 55827 30685
rect 55861 30719 55919 30725
rect 55861 30685 55873 30719
rect 55907 30685 55919 30719
rect 57146 30716 57152 30728
rect 57107 30688 57152 30716
rect 55861 30679 55919 30685
rect 50672 30620 51304 30648
rect 51353 30651 51411 30657
rect 50672 30608 50678 30620
rect 51353 30617 51365 30651
rect 51399 30648 51411 30651
rect 51994 30648 52000 30660
rect 51399 30620 52000 30648
rect 51399 30617 51411 30620
rect 51353 30611 51411 30617
rect 51994 30608 52000 30620
rect 52052 30608 52058 30660
rect 52178 30608 52184 30660
rect 52236 30648 52242 30660
rect 52822 30648 52828 30660
rect 52236 30620 52684 30648
rect 52783 30620 52828 30648
rect 52236 30608 52242 30620
rect 47728 30552 47809 30580
rect 52273 30583 52331 30589
rect 47728 30540 47734 30552
rect 52273 30549 52285 30583
rect 52319 30580 52331 30583
rect 52362 30580 52368 30592
rect 52319 30552 52368 30580
rect 52319 30549 52331 30552
rect 52273 30543 52331 30549
rect 52362 30540 52368 30552
rect 52420 30540 52426 30592
rect 52656 30580 52684 30620
rect 52822 30608 52828 30620
rect 52880 30608 52886 30660
rect 52917 30651 52975 30657
rect 52917 30617 52929 30651
rect 52963 30648 52975 30651
rect 54110 30648 54116 30660
rect 52963 30620 54116 30648
rect 52963 30617 52975 30620
rect 52917 30611 52975 30617
rect 52932 30580 52960 30611
rect 54110 30608 54116 30620
rect 54168 30608 54174 30660
rect 54570 30648 54576 30660
rect 54531 30620 54576 30648
rect 54570 30608 54576 30620
rect 54628 30608 54634 30660
rect 54665 30651 54723 30657
rect 54665 30617 54677 30651
rect 54711 30617 54723 30651
rect 54665 30611 54723 30617
rect 52656 30552 52960 30580
rect 53834 30540 53840 30592
rect 53892 30580 53898 30592
rect 54021 30583 54079 30589
rect 54021 30580 54033 30583
rect 53892 30552 54033 30580
rect 53892 30540 53898 30552
rect 54021 30549 54033 30552
rect 54067 30549 54079 30583
rect 54128 30580 54156 30608
rect 54680 30580 54708 30611
rect 54938 30608 54944 30660
rect 54996 30648 55002 30660
rect 55876 30648 55904 30679
rect 57146 30676 57152 30688
rect 57204 30676 57210 30728
rect 54996 30620 55904 30648
rect 54996 30608 55002 30620
rect 56502 30608 56508 30660
rect 56560 30648 56566 30660
rect 57977 30651 58035 30657
rect 57977 30648 57989 30651
rect 56560 30620 57989 30648
rect 56560 30608 56566 30620
rect 57977 30617 57989 30620
rect 58023 30617 58035 30651
rect 57977 30611 58035 30617
rect 54128 30552 54708 30580
rect 56045 30583 56103 30589
rect 54021 30543 54079 30549
rect 56045 30549 56057 30583
rect 56091 30580 56103 30583
rect 57054 30580 57060 30592
rect 56091 30552 57060 30580
rect 56091 30549 56103 30552
rect 56045 30543 56103 30549
rect 57054 30540 57060 30552
rect 57112 30540 57118 30592
rect 1104 30490 58880 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 58880 30490
rect 1104 30416 58880 30438
rect 34698 30336 34704 30388
rect 34756 30336 34762 30388
rect 34790 30336 34796 30388
rect 34848 30376 34854 30388
rect 34848 30348 34928 30376
rect 34848 30336 34854 30348
rect 30834 30308 30840 30320
rect 30795 30280 30840 30308
rect 30834 30268 30840 30280
rect 30892 30268 30898 30320
rect 33873 30311 33931 30317
rect 33873 30277 33885 30311
rect 33919 30308 33931 30311
rect 34716 30308 34744 30336
rect 34900 30317 34928 30348
rect 35158 30336 35164 30388
rect 35216 30376 35222 30388
rect 35618 30376 35624 30388
rect 35216 30348 35624 30376
rect 35216 30336 35222 30348
rect 35618 30336 35624 30348
rect 35676 30336 35682 30388
rect 36354 30376 36360 30388
rect 36315 30348 36360 30376
rect 36354 30336 36360 30348
rect 36412 30336 36418 30388
rect 36722 30336 36728 30388
rect 36780 30376 36786 30388
rect 37274 30376 37280 30388
rect 36780 30348 37280 30376
rect 36780 30336 36786 30348
rect 37274 30336 37280 30348
rect 37332 30376 37338 30388
rect 41046 30376 41052 30388
rect 37332 30348 37780 30376
rect 37332 30336 37338 30348
rect 33919 30280 34744 30308
rect 34885 30311 34943 30317
rect 33919 30277 33931 30280
rect 33873 30271 33931 30277
rect 34885 30277 34897 30311
rect 34931 30277 34943 30311
rect 34885 30271 34943 30277
rect 35342 30268 35348 30320
rect 35400 30268 35406 30320
rect 37550 30268 37556 30320
rect 37608 30268 37614 30320
rect 37752 30317 37780 30348
rect 40282 30348 41052 30376
rect 37737 30311 37795 30317
rect 37737 30277 37749 30311
rect 37783 30277 37795 30311
rect 37737 30271 37795 30277
rect 37918 30268 37924 30320
rect 37976 30317 37982 30320
rect 37976 30311 38005 30317
rect 37993 30277 38005 30311
rect 37976 30271 38005 30277
rect 37976 30268 37982 30271
rect 38562 30268 38568 30320
rect 38620 30308 38626 30320
rect 38620 30280 39988 30308
rect 38620 30268 38626 30280
rect 28810 30240 28816 30252
rect 28771 30212 28816 30240
rect 28810 30200 28816 30212
rect 28868 30200 28874 30252
rect 28902 30200 28908 30252
rect 28960 30240 28966 30252
rect 29457 30243 29515 30249
rect 29457 30240 29469 30243
rect 28960 30212 29469 30240
rect 28960 30200 28966 30212
rect 29457 30209 29469 30212
rect 29503 30240 29515 30243
rect 29917 30243 29975 30249
rect 29917 30240 29929 30243
rect 29503 30212 29929 30240
rect 29503 30209 29515 30212
rect 29457 30203 29515 30209
rect 29917 30209 29929 30212
rect 29963 30209 29975 30243
rect 29917 30203 29975 30209
rect 29932 30172 29960 30203
rect 30282 30200 30288 30252
rect 30340 30240 30346 30252
rect 30929 30243 30987 30249
rect 30929 30240 30941 30243
rect 30340 30212 30941 30240
rect 30340 30200 30346 30212
rect 30929 30209 30941 30212
rect 30975 30240 30987 30243
rect 31754 30240 31760 30252
rect 30975 30212 31760 30240
rect 30975 30209 30987 30212
rect 30929 30203 30987 30209
rect 31754 30200 31760 30212
rect 31812 30200 31818 30252
rect 32766 30200 32772 30252
rect 32824 30200 32830 30252
rect 34146 30200 34152 30252
rect 34204 30240 34210 30252
rect 34609 30243 34667 30249
rect 34609 30240 34621 30243
rect 34204 30212 34621 30240
rect 34204 30200 34210 30212
rect 34609 30209 34621 30212
rect 34655 30209 34667 30243
rect 37568 30240 37596 30268
rect 39960 30252 39988 30280
rect 40034 30268 40040 30320
rect 40092 30308 40098 30320
rect 40282 30317 40310 30348
rect 41046 30336 41052 30348
rect 41104 30336 41110 30388
rect 47670 30376 47676 30388
rect 46492 30348 47676 30376
rect 40267 30311 40325 30317
rect 40092 30280 40137 30308
rect 40092 30268 40098 30280
rect 40267 30277 40279 30311
rect 40313 30277 40325 30311
rect 40678 30308 40684 30320
rect 40267 30271 40325 30277
rect 40420 30280 40684 30308
rect 37645 30243 37703 30249
rect 37645 30240 37657 30243
rect 37568 30212 37657 30240
rect 34609 30203 34667 30209
rect 37645 30209 37657 30212
rect 37691 30209 37703 30243
rect 37645 30203 37703 30209
rect 37826 30200 37832 30252
rect 37884 30240 37890 30252
rect 37884 30212 37964 30240
rect 37884 30200 37890 30212
rect 29932 30144 34744 30172
rect 28534 30064 28540 30116
rect 28592 30104 28598 30116
rect 28629 30107 28687 30113
rect 28629 30104 28641 30107
rect 28592 30076 28641 30104
rect 28592 30064 28598 30076
rect 28629 30073 28641 30076
rect 28675 30073 28687 30107
rect 28629 30067 28687 30073
rect 30101 30107 30159 30113
rect 30101 30073 30113 30107
rect 30147 30104 30159 30107
rect 30147 30076 32904 30104
rect 30147 30073 30159 30076
rect 30101 30067 30159 30073
rect 31481 30039 31539 30045
rect 31481 30005 31493 30039
rect 31527 30036 31539 30039
rect 31754 30036 31760 30048
rect 31527 30008 31760 30036
rect 31527 30005 31539 30008
rect 31481 29999 31539 30005
rect 31754 29996 31760 30008
rect 31812 29996 31818 30048
rect 32398 30036 32404 30048
rect 32359 30008 32404 30036
rect 32398 29996 32404 30008
rect 32456 29996 32462 30048
rect 32876 30036 32904 30076
rect 34716 30048 34744 30144
rect 34882 30132 34888 30184
rect 34940 30172 34946 30184
rect 37461 30175 37519 30181
rect 37461 30172 37473 30175
rect 34940 30144 37473 30172
rect 34940 30132 34946 30144
rect 37461 30141 37473 30144
rect 37507 30141 37519 30175
rect 37936 30172 37964 30212
rect 38102 30200 38108 30252
rect 38160 30240 38166 30252
rect 38160 30212 38205 30240
rect 38160 30200 38166 30212
rect 38654 30200 38660 30252
rect 38712 30240 38718 30252
rect 38749 30243 38807 30249
rect 38749 30240 38761 30243
rect 38712 30212 38761 30240
rect 38712 30200 38718 30212
rect 38749 30209 38761 30212
rect 38795 30209 38807 30243
rect 39942 30240 39948 30252
rect 38749 30203 38807 30209
rect 38856 30212 39160 30240
rect 39903 30212 39948 30240
rect 38856 30172 38884 30212
rect 37936 30144 38884 30172
rect 38933 30175 38991 30181
rect 37461 30135 37519 30141
rect 38933 30141 38945 30175
rect 38979 30172 38991 30175
rect 39022 30172 39028 30184
rect 38979 30144 39028 30172
rect 38979 30141 38991 30144
rect 38933 30135 38991 30141
rect 39022 30132 39028 30144
rect 39080 30132 39086 30184
rect 39132 30172 39160 30212
rect 39942 30200 39948 30212
rect 40000 30200 40006 30252
rect 40129 30243 40187 30249
rect 40129 30209 40141 30243
rect 40175 30209 40187 30243
rect 40129 30203 40187 30209
rect 39206 30172 39212 30184
rect 39132 30144 39212 30172
rect 39206 30132 39212 30144
rect 39264 30172 39270 30184
rect 40144 30172 40172 30203
rect 40420 30184 40448 30280
rect 40678 30268 40684 30280
rect 40736 30268 40742 30320
rect 40862 30268 40868 30320
rect 40920 30308 40926 30320
rect 41325 30311 41383 30317
rect 41325 30308 41337 30311
rect 40920 30280 41337 30308
rect 40920 30268 40926 30280
rect 41325 30277 41337 30280
rect 41371 30277 41383 30311
rect 45186 30308 45192 30320
rect 45147 30280 45192 30308
rect 41325 30271 41383 30277
rect 45186 30268 45192 30280
rect 45244 30268 45250 30320
rect 45738 30268 45744 30320
rect 45796 30308 45802 30320
rect 46492 30308 46520 30348
rect 47670 30336 47676 30348
rect 47728 30336 47734 30388
rect 47857 30379 47915 30385
rect 47857 30345 47869 30379
rect 47903 30376 47915 30379
rect 48314 30376 48320 30388
rect 47903 30348 48320 30376
rect 47903 30345 47915 30348
rect 47857 30339 47915 30345
rect 48314 30336 48320 30348
rect 48372 30376 48378 30388
rect 51166 30376 51172 30388
rect 48372 30348 51172 30376
rect 48372 30336 48378 30348
rect 48501 30311 48559 30317
rect 48501 30308 48513 30311
rect 45796 30280 46520 30308
rect 45796 30268 45802 30280
rect 40494 30200 40500 30252
rect 40552 30240 40558 30252
rect 41187 30243 41245 30249
rect 41187 30240 41199 30243
rect 40552 30212 41199 30240
rect 40552 30200 40558 30212
rect 41187 30209 41199 30212
rect 41233 30209 41245 30243
rect 41416 30243 41474 30249
rect 41416 30240 41428 30243
rect 41187 30203 41245 30209
rect 41340 30212 41428 30240
rect 41340 30184 41368 30212
rect 41416 30209 41428 30212
rect 41462 30209 41474 30243
rect 41416 30203 41474 30209
rect 41506 30200 41512 30252
rect 41564 30240 41570 30252
rect 41564 30212 41608 30240
rect 41564 30200 41570 30212
rect 42794 30200 42800 30252
rect 42852 30240 42858 30252
rect 43162 30240 43168 30252
rect 42852 30212 43168 30240
rect 42852 30200 42858 30212
rect 43162 30200 43168 30212
rect 43220 30200 43226 30252
rect 44542 30200 44548 30252
rect 44600 30200 44606 30252
rect 45554 30200 45560 30252
rect 45612 30240 45618 30252
rect 46293 30243 46351 30249
rect 46293 30240 46305 30243
rect 45612 30212 46305 30240
rect 45612 30200 45618 30212
rect 46293 30209 46305 30212
rect 46339 30209 46351 30243
rect 46293 30203 46351 30209
rect 46385 30243 46443 30249
rect 46385 30209 46397 30243
rect 46431 30240 46443 30243
rect 46492 30240 46520 30280
rect 46584 30280 48513 30308
rect 46584 30249 46612 30280
rect 48501 30277 48513 30280
rect 48547 30277 48559 30311
rect 49694 30308 49700 30320
rect 49607 30280 49700 30308
rect 48501 30271 48559 30277
rect 49694 30268 49700 30280
rect 49752 30308 49758 30320
rect 50430 30308 50436 30320
rect 49752 30280 50436 30308
rect 49752 30268 49758 30280
rect 50430 30268 50436 30280
rect 50488 30268 50494 30320
rect 46431 30212 46520 30240
rect 46569 30243 46627 30249
rect 46431 30209 46443 30212
rect 46385 30203 46443 30209
rect 46569 30209 46581 30243
rect 46615 30209 46627 30243
rect 46569 30203 46627 30209
rect 46658 30200 46664 30252
rect 46716 30240 46722 30252
rect 46716 30212 46761 30240
rect 46716 30200 46722 30212
rect 46842 30200 46848 30252
rect 46900 30240 46906 30252
rect 47121 30243 47179 30249
rect 47121 30240 47133 30243
rect 46900 30212 47133 30240
rect 46900 30200 46906 30212
rect 47121 30209 47133 30212
rect 47167 30209 47179 30243
rect 47121 30203 47179 30209
rect 47765 30243 47823 30249
rect 47765 30209 47777 30243
rect 47811 30209 47823 30243
rect 47765 30203 47823 30209
rect 47949 30243 48007 30249
rect 47949 30209 47961 30243
rect 47995 30240 48007 30243
rect 48314 30240 48320 30252
rect 47995 30212 48320 30240
rect 47995 30209 48007 30212
rect 47949 30203 48007 30209
rect 40402 30172 40408 30184
rect 39264 30144 40172 30172
rect 40363 30144 40408 30172
rect 39264 30132 39270 30144
rect 35894 30064 35900 30116
rect 35952 30104 35958 30116
rect 39761 30107 39819 30113
rect 39761 30104 39773 30107
rect 35952 30076 39773 30104
rect 35952 30064 35958 30076
rect 39761 30073 39773 30076
rect 39807 30073 39819 30107
rect 40144 30104 40172 30144
rect 40402 30132 40408 30144
rect 40460 30132 40466 30184
rect 41049 30175 41107 30181
rect 41049 30141 41061 30175
rect 41095 30141 41107 30175
rect 41049 30135 41107 30141
rect 40310 30104 40316 30116
rect 40144 30076 40316 30104
rect 39761 30067 39819 30073
rect 40310 30064 40316 30076
rect 40368 30104 40374 30116
rect 40678 30104 40684 30116
rect 40368 30076 40684 30104
rect 40368 30064 40374 30076
rect 40678 30064 40684 30076
rect 40736 30104 40742 30116
rect 40862 30104 40868 30116
rect 40736 30076 40868 30104
rect 40736 30064 40742 30076
rect 40862 30064 40868 30076
rect 40920 30064 40926 30116
rect 41064 30104 41092 30135
rect 41322 30132 41328 30184
rect 41380 30132 41386 30184
rect 41693 30175 41751 30181
rect 41693 30141 41705 30175
rect 41739 30172 41751 30175
rect 43441 30175 43499 30181
rect 43441 30172 43453 30175
rect 41739 30144 43453 30172
rect 41739 30141 41751 30144
rect 41693 30135 41751 30141
rect 43441 30141 43453 30144
rect 43487 30141 43499 30175
rect 43441 30135 43499 30141
rect 45278 30132 45284 30184
rect 45336 30172 45342 30184
rect 47670 30172 47676 30184
rect 45336 30144 47676 30172
rect 45336 30132 45342 30144
rect 47670 30132 47676 30144
rect 47728 30172 47734 30184
rect 47780 30172 47808 30203
rect 48314 30200 48320 30212
rect 48372 30200 48378 30252
rect 48409 30243 48467 30249
rect 48409 30209 48421 30243
rect 48455 30209 48467 30243
rect 48409 30203 48467 30209
rect 48593 30243 48651 30249
rect 48593 30209 48605 30243
rect 48639 30240 48651 30243
rect 48866 30240 48872 30252
rect 48639 30212 48872 30240
rect 48639 30209 48651 30212
rect 48593 30203 48651 30209
rect 47728 30144 47808 30172
rect 47728 30132 47734 30144
rect 42978 30104 42984 30116
rect 41064 30076 42984 30104
rect 42978 30064 42984 30076
rect 43036 30064 43042 30116
rect 46290 30064 46296 30116
rect 46348 30104 46354 30116
rect 48424 30104 48452 30203
rect 48866 30200 48872 30212
rect 48924 30200 48930 30252
rect 50540 30249 50568 30348
rect 51166 30336 51172 30348
rect 51224 30336 51230 30388
rect 52178 30336 52184 30388
rect 52236 30336 52242 30388
rect 53374 30376 53380 30388
rect 52288 30348 53380 30376
rect 50614 30268 50620 30320
rect 50672 30308 50678 30320
rect 50985 30311 51043 30317
rect 50672 30280 50717 30308
rect 50672 30268 50678 30280
rect 50985 30277 50997 30311
rect 51031 30308 51043 30311
rect 52196 30308 52224 30336
rect 51031 30280 52224 30308
rect 51031 30277 51043 30280
rect 50985 30271 51043 30277
rect 49329 30243 49387 30249
rect 49329 30240 49341 30243
rect 48976 30212 49341 30240
rect 48498 30132 48504 30184
rect 48556 30172 48562 30184
rect 48976 30172 49004 30212
rect 49329 30209 49341 30212
rect 49375 30209 49387 30243
rect 49329 30203 49387 30209
rect 50525 30243 50583 30249
rect 50525 30209 50537 30243
rect 50571 30209 50583 30243
rect 50798 30240 50804 30252
rect 50759 30212 50804 30240
rect 50525 30203 50583 30209
rect 50798 30200 50804 30212
rect 50856 30200 50862 30252
rect 51994 30240 52000 30252
rect 51907 30212 52000 30240
rect 51994 30200 52000 30212
rect 52052 30200 52058 30252
rect 52089 30243 52147 30249
rect 52089 30209 52101 30243
rect 52135 30240 52147 30243
rect 52178 30240 52184 30252
rect 52135 30212 52184 30240
rect 52135 30209 52147 30212
rect 52089 30203 52147 30209
rect 52178 30200 52184 30212
rect 52236 30200 52242 30252
rect 52288 30249 52316 30348
rect 53374 30336 53380 30348
rect 53432 30336 53438 30388
rect 53581 30348 54064 30376
rect 52273 30243 52331 30249
rect 52273 30209 52285 30243
rect 52319 30209 52331 30243
rect 52273 30203 52331 30209
rect 52362 30200 52368 30252
rect 52420 30240 52426 30252
rect 53193 30243 53251 30249
rect 52420 30212 52465 30240
rect 52420 30200 52426 30212
rect 53193 30209 53205 30243
rect 53239 30240 53251 30243
rect 53581 30240 53609 30348
rect 53834 30308 53840 30320
rect 53668 30280 53840 30308
rect 53668 30249 53696 30280
rect 53834 30268 53840 30280
rect 53892 30268 53898 30320
rect 53239 30212 53609 30240
rect 53653 30243 53711 30249
rect 53239 30209 53251 30212
rect 53193 30203 53251 30209
rect 53653 30209 53665 30243
rect 53699 30209 53711 30243
rect 53653 30203 53711 30209
rect 48556 30144 49004 30172
rect 48556 30132 48562 30144
rect 49142 30132 49148 30184
rect 49200 30172 49206 30184
rect 52012 30172 52040 30200
rect 53208 30172 53236 30203
rect 53742 30200 53748 30252
rect 53800 30240 53806 30252
rect 53926 30240 53932 30252
rect 53800 30212 53845 30240
rect 53887 30212 53932 30240
rect 53800 30200 53806 30212
rect 53926 30200 53932 30212
rect 53984 30200 53990 30252
rect 54036 30249 54064 30348
rect 54110 30336 54116 30388
rect 54168 30376 54174 30388
rect 54168 30348 55352 30376
rect 54168 30336 54174 30348
rect 55324 30320 55352 30348
rect 57882 30336 57888 30388
rect 57940 30376 57946 30388
rect 57940 30348 58112 30376
rect 57940 30336 57946 30348
rect 54757 30311 54815 30317
rect 54757 30277 54769 30311
rect 54803 30308 54815 30311
rect 55030 30308 55036 30320
rect 54803 30280 55036 30308
rect 54803 30277 54815 30280
rect 54757 30271 54815 30277
rect 55030 30268 55036 30280
rect 55088 30268 55094 30320
rect 55306 30268 55312 30320
rect 55364 30308 55370 30320
rect 56321 30311 56379 30317
rect 56321 30308 56333 30311
rect 55364 30280 56333 30308
rect 55364 30268 55370 30280
rect 56321 30277 56333 30280
rect 56367 30308 56379 30311
rect 56594 30308 56600 30320
rect 56367 30280 56600 30308
rect 56367 30277 56379 30280
rect 56321 30271 56379 30277
rect 56594 30268 56600 30280
rect 56652 30268 56658 30320
rect 58084 30317 58112 30348
rect 58069 30311 58127 30317
rect 58069 30277 58081 30311
rect 58115 30277 58127 30311
rect 58069 30271 58127 30277
rect 54021 30243 54079 30249
rect 54021 30209 54033 30243
rect 54067 30240 54079 30243
rect 54202 30240 54208 30252
rect 54067 30212 54208 30240
rect 54067 30209 54079 30212
rect 54021 30203 54079 30209
rect 54202 30200 54208 30212
rect 54260 30240 54266 30252
rect 54938 30240 54944 30252
rect 54260 30212 54944 30240
rect 54260 30200 54266 30212
rect 54938 30200 54944 30212
rect 54996 30200 55002 30252
rect 55766 30200 55772 30252
rect 55824 30240 55830 30252
rect 56045 30243 56103 30249
rect 56045 30240 56057 30243
rect 55824 30212 56057 30240
rect 55824 30200 55830 30212
rect 56045 30209 56057 30212
rect 56091 30240 56103 30243
rect 56134 30240 56140 30252
rect 56091 30212 56140 30240
rect 56091 30209 56103 30212
rect 56045 30203 56103 30209
rect 56134 30200 56140 30212
rect 56192 30200 56198 30252
rect 57149 30243 57207 30249
rect 57149 30209 57161 30243
rect 57195 30240 57207 30243
rect 57330 30240 57336 30252
rect 57195 30212 57336 30240
rect 57195 30209 57207 30212
rect 57149 30203 57207 30209
rect 57330 30200 57336 30212
rect 57388 30200 57394 30252
rect 49200 30144 49245 30172
rect 52012 30144 53236 30172
rect 49200 30132 49206 30144
rect 53282 30132 53288 30184
rect 53340 30172 53346 30184
rect 55217 30175 55275 30181
rect 55217 30172 55229 30175
rect 53340 30144 55229 30172
rect 53340 30132 53346 30144
rect 55217 30141 55229 30144
rect 55263 30141 55275 30175
rect 55217 30135 55275 30141
rect 55490 30132 55496 30184
rect 55548 30172 55554 30184
rect 55953 30175 56011 30181
rect 55953 30172 55965 30175
rect 55548 30144 55965 30172
rect 55548 30132 55554 30144
rect 55953 30141 55965 30144
rect 55999 30141 56011 30175
rect 56410 30172 56416 30184
rect 56371 30144 56416 30172
rect 55953 30135 56011 30141
rect 46348 30076 48452 30104
rect 49605 30107 49663 30113
rect 46348 30064 46354 30076
rect 49605 30073 49617 30107
rect 49651 30104 49663 30107
rect 52546 30104 52552 30116
rect 49651 30076 52552 30104
rect 49651 30073 49663 30076
rect 49605 30067 49663 30073
rect 52546 30064 52552 30076
rect 52604 30064 52610 30116
rect 55968 30104 55996 30135
rect 56410 30132 56416 30144
rect 56468 30132 56474 30184
rect 57054 30172 57060 30184
rect 57015 30144 57060 30172
rect 57054 30132 57060 30144
rect 57112 30132 57118 30184
rect 56042 30104 56048 30116
rect 55968 30076 56048 30104
rect 56042 30064 56048 30076
rect 56100 30064 56106 30116
rect 57514 30104 57520 30116
rect 57475 30076 57520 30104
rect 57514 30064 57520 30076
rect 57572 30064 57578 30116
rect 34514 30036 34520 30048
rect 32876 30008 34520 30036
rect 34514 29996 34520 30008
rect 34572 29996 34578 30048
rect 34698 29996 34704 30048
rect 34756 30036 34762 30048
rect 35434 30036 35440 30048
rect 34756 30008 35440 30036
rect 34756 29996 34762 30008
rect 35434 29996 35440 30008
rect 35492 29996 35498 30048
rect 35526 29996 35532 30048
rect 35584 30036 35590 30048
rect 38194 30036 38200 30048
rect 35584 30008 38200 30036
rect 35584 29996 35590 30008
rect 38194 29996 38200 30008
rect 38252 29996 38258 30048
rect 38470 29996 38476 30048
rect 38528 30036 38534 30048
rect 38565 30039 38623 30045
rect 38565 30036 38577 30039
rect 38528 30008 38577 30036
rect 38528 29996 38534 30008
rect 38565 30005 38577 30008
rect 38611 30036 38623 30039
rect 41506 30036 41512 30048
rect 38611 30008 41512 30036
rect 38611 30005 38623 30008
rect 38565 29999 38623 30005
rect 41506 29996 41512 30008
rect 41564 29996 41570 30048
rect 41598 29996 41604 30048
rect 41656 30036 41662 30048
rect 42613 30039 42671 30045
rect 42613 30036 42625 30039
rect 41656 30008 42625 30036
rect 41656 29996 41662 30008
rect 42613 30005 42625 30008
rect 42659 30005 42671 30039
rect 42613 29999 42671 30005
rect 46109 30039 46167 30045
rect 46109 30005 46121 30039
rect 46155 30036 46167 30039
rect 50246 30036 50252 30048
rect 46155 30008 50252 30036
rect 46155 30005 46167 30008
rect 46109 29999 46167 30005
rect 50246 29996 50252 30008
rect 50304 29996 50310 30048
rect 51813 30039 51871 30045
rect 51813 30005 51825 30039
rect 51859 30036 51871 30039
rect 51902 30036 51908 30048
rect 51859 30008 51908 30036
rect 51859 30005 51871 30008
rect 51813 29999 51871 30005
rect 51902 29996 51908 30008
rect 51960 29996 51966 30048
rect 53009 30039 53067 30045
rect 53009 30005 53021 30039
rect 53055 30036 53067 30039
rect 53098 30036 53104 30048
rect 53055 30008 53104 30036
rect 53055 30005 53067 30008
rect 53009 29999 53067 30005
rect 53098 29996 53104 30008
rect 53156 30036 53162 30048
rect 53558 30036 53564 30048
rect 53156 30008 53564 30036
rect 53156 29996 53162 30008
rect 53558 29996 53564 30008
rect 53616 29996 53622 30048
rect 54205 30039 54263 30045
rect 54205 30005 54217 30039
rect 54251 30036 54263 30039
rect 55122 30036 55128 30048
rect 54251 30008 55128 30036
rect 54251 30005 54263 30008
rect 54205 29999 54263 30005
rect 55122 29996 55128 30008
rect 55180 29996 55186 30048
rect 55769 30039 55827 30045
rect 55769 30005 55781 30039
rect 55815 30036 55827 30039
rect 55950 30036 55956 30048
rect 55815 30008 55956 30036
rect 55815 30005 55827 30008
rect 55769 29999 55827 30005
rect 55950 29996 55956 30008
rect 56008 29996 56014 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 29362 29792 29368 29844
rect 29420 29832 29426 29844
rect 29825 29835 29883 29841
rect 29825 29832 29837 29835
rect 29420 29804 29837 29832
rect 29420 29792 29426 29804
rect 29825 29801 29837 29804
rect 29871 29801 29883 29835
rect 29825 29795 29883 29801
rect 31846 29792 31852 29844
rect 31904 29832 31910 29844
rect 32493 29835 32551 29841
rect 32493 29832 32505 29835
rect 31904 29804 32505 29832
rect 31904 29792 31910 29804
rect 32493 29801 32505 29804
rect 32539 29832 32551 29835
rect 33410 29832 33416 29844
rect 32539 29804 33416 29832
rect 32539 29801 32551 29804
rect 32493 29795 32551 29801
rect 33410 29792 33416 29804
rect 33468 29832 33474 29844
rect 34146 29832 34152 29844
rect 33468 29804 34152 29832
rect 33468 29792 33474 29804
rect 34146 29792 34152 29804
rect 34204 29792 34210 29844
rect 34977 29835 35035 29841
rect 34977 29801 34989 29835
rect 35023 29832 35035 29835
rect 35342 29832 35348 29844
rect 35023 29804 35348 29832
rect 35023 29801 35035 29804
rect 34977 29795 35035 29801
rect 35342 29792 35348 29804
rect 35400 29792 35406 29844
rect 36446 29832 36452 29844
rect 36407 29804 36452 29832
rect 36446 29792 36452 29804
rect 36504 29792 36510 29844
rect 40773 29835 40831 29841
rect 40773 29832 40785 29835
rect 36556 29804 40785 29832
rect 31573 29699 31631 29705
rect 31573 29665 31585 29699
rect 31619 29696 31631 29699
rect 31864 29696 31892 29792
rect 35894 29764 35900 29776
rect 31619 29668 31892 29696
rect 34072 29736 35900 29764
rect 31619 29665 31631 29668
rect 31573 29659 31631 29665
rect 30190 29588 30196 29640
rect 30248 29588 30254 29640
rect 31662 29588 31668 29640
rect 31720 29628 31726 29640
rect 34072 29628 34100 29736
rect 35894 29724 35900 29736
rect 35952 29724 35958 29776
rect 36556 29696 36584 29804
rect 40773 29801 40785 29804
rect 40819 29801 40831 29835
rect 41782 29832 41788 29844
rect 40773 29795 40831 29801
rect 41222 29804 41788 29832
rect 37550 29764 37556 29776
rect 31720 29600 34100 29628
rect 34256 29668 36584 29696
rect 36648 29736 37556 29764
rect 31720 29588 31726 29600
rect 31294 29560 31300 29572
rect 31255 29532 31300 29560
rect 31294 29520 31300 29532
rect 31352 29520 31358 29572
rect 32950 29520 32956 29572
rect 33008 29560 33014 29572
rect 33781 29563 33839 29569
rect 33781 29560 33793 29563
rect 33008 29532 33793 29560
rect 33008 29520 33014 29532
rect 33781 29529 33793 29532
rect 33827 29529 33839 29563
rect 33781 29523 33839 29529
rect 28810 29452 28816 29504
rect 28868 29492 28874 29504
rect 34256 29492 34284 29668
rect 34790 29588 34796 29640
rect 34848 29628 34854 29640
rect 34885 29631 34943 29637
rect 34885 29628 34897 29631
rect 34848 29600 34897 29628
rect 34848 29588 34854 29600
rect 34885 29597 34897 29600
rect 34931 29628 34943 29631
rect 35526 29628 35532 29640
rect 34931 29600 35532 29628
rect 34931 29597 34943 29600
rect 34885 29591 34943 29597
rect 35526 29588 35532 29600
rect 35584 29588 35590 29640
rect 36648 29637 36676 29736
rect 37550 29724 37556 29736
rect 37608 29764 37614 29776
rect 38562 29764 38568 29776
rect 37608 29736 38568 29764
rect 37608 29724 37614 29736
rect 38562 29724 38568 29736
rect 38620 29724 38626 29776
rect 38657 29767 38715 29773
rect 38657 29733 38669 29767
rect 38703 29764 38715 29767
rect 39758 29764 39764 29776
rect 38703 29736 39764 29764
rect 38703 29733 38715 29736
rect 38657 29727 38715 29733
rect 39758 29724 39764 29736
rect 39816 29724 39822 29776
rect 40126 29724 40132 29776
rect 40184 29764 40190 29776
rect 40402 29764 40408 29776
rect 40184 29736 40408 29764
rect 40184 29724 40190 29736
rect 40402 29724 40408 29736
rect 40460 29724 40466 29776
rect 37093 29699 37151 29705
rect 37093 29665 37105 29699
rect 37139 29696 37151 29699
rect 37366 29696 37372 29708
rect 37139 29668 37372 29696
rect 37139 29665 37151 29668
rect 37093 29659 37151 29665
rect 37366 29656 37372 29668
rect 37424 29656 37430 29708
rect 37921 29699 37979 29705
rect 37921 29665 37933 29699
rect 37967 29696 37979 29699
rect 38930 29696 38936 29708
rect 37967 29668 38936 29696
rect 37967 29665 37979 29668
rect 37921 29659 37979 29665
rect 38930 29656 38936 29668
rect 38988 29696 38994 29708
rect 41222 29705 41250 29804
rect 41782 29792 41788 29804
rect 41840 29832 41846 29844
rect 42702 29832 42708 29844
rect 41840 29804 42708 29832
rect 41840 29792 41846 29804
rect 42702 29792 42708 29804
rect 42760 29792 42766 29844
rect 44542 29832 44548 29844
rect 44503 29804 44548 29832
rect 44542 29792 44548 29804
rect 44600 29792 44606 29844
rect 46382 29832 46388 29844
rect 46343 29804 46388 29832
rect 46382 29792 46388 29804
rect 46440 29792 46446 29844
rect 46477 29835 46535 29841
rect 46477 29801 46489 29835
rect 46523 29832 46535 29835
rect 46658 29832 46664 29844
rect 46523 29804 46664 29832
rect 46523 29801 46535 29804
rect 46477 29795 46535 29801
rect 46658 29792 46664 29804
rect 46716 29792 46722 29844
rect 47210 29832 47216 29844
rect 47171 29804 47216 29832
rect 47210 29792 47216 29804
rect 47268 29792 47274 29844
rect 47670 29792 47676 29844
rect 47728 29832 47734 29844
rect 49142 29832 49148 29844
rect 47728 29804 49148 29832
rect 47728 29792 47734 29804
rect 49142 29792 49148 29804
rect 49200 29832 49206 29844
rect 49237 29835 49295 29841
rect 49237 29832 49249 29835
rect 49200 29804 49249 29832
rect 49200 29792 49206 29804
rect 49237 29801 49249 29804
rect 49283 29801 49295 29835
rect 49237 29795 49295 29801
rect 49421 29835 49479 29841
rect 49421 29801 49433 29835
rect 49467 29832 49479 29835
rect 53742 29832 53748 29844
rect 49467 29804 53748 29832
rect 49467 29801 49479 29804
rect 49421 29795 49479 29801
rect 53742 29792 53748 29804
rect 53800 29792 53806 29844
rect 41322 29724 41328 29776
rect 41380 29764 41386 29776
rect 45833 29767 45891 29773
rect 41380 29736 41459 29764
rect 41380 29724 41386 29736
rect 41431 29705 41459 29736
rect 45833 29733 45845 29767
rect 45879 29764 45891 29767
rect 47578 29764 47584 29776
rect 45879 29736 47584 29764
rect 45879 29733 45891 29736
rect 45833 29727 45891 29733
rect 47578 29724 47584 29736
rect 47636 29724 47642 29776
rect 47857 29767 47915 29773
rect 47857 29733 47869 29767
rect 47903 29764 47915 29767
rect 49050 29764 49056 29776
rect 47903 29736 49056 29764
rect 47903 29733 47915 29736
rect 47857 29727 47915 29733
rect 49050 29724 49056 29736
rect 49108 29724 49114 29776
rect 56502 29764 56508 29776
rect 54128 29736 56508 29764
rect 39025 29699 39083 29705
rect 39025 29696 39037 29699
rect 38988 29668 39037 29696
rect 38988 29656 38994 29668
rect 39025 29665 39037 29668
rect 39071 29696 39083 29699
rect 41222 29699 41291 29705
rect 41222 29696 41245 29699
rect 39071 29668 41245 29696
rect 39071 29665 39083 29668
rect 39025 29659 39083 29665
rect 41233 29665 41245 29668
rect 41279 29665 41291 29699
rect 41233 29659 41291 29665
rect 41417 29699 41475 29705
rect 41417 29665 41429 29699
rect 41463 29665 41475 29699
rect 41417 29659 41475 29665
rect 41969 29699 42027 29705
rect 41969 29665 41981 29699
rect 42015 29696 42027 29699
rect 42794 29696 42800 29708
rect 42015 29668 42800 29696
rect 42015 29665 42027 29668
rect 41969 29659 42027 29665
rect 42794 29656 42800 29668
rect 42852 29656 42858 29708
rect 44266 29656 44272 29708
rect 44324 29696 44330 29708
rect 44324 29668 45508 29696
rect 44324 29656 44330 29668
rect 36633 29631 36691 29637
rect 36633 29597 36645 29631
rect 36679 29597 36691 29631
rect 36814 29628 36820 29640
rect 36775 29600 36820 29628
rect 36633 29591 36691 29597
rect 36814 29588 36820 29600
rect 36872 29588 36878 29640
rect 37737 29631 37795 29637
rect 37737 29597 37749 29631
rect 37783 29597 37795 29631
rect 37737 29591 37795 29597
rect 34330 29520 34336 29572
rect 34388 29560 34394 29572
rect 35986 29560 35992 29572
rect 34388 29532 35992 29560
rect 34388 29520 34394 29532
rect 35986 29520 35992 29532
rect 36044 29520 36050 29572
rect 36725 29563 36783 29569
rect 36725 29529 36737 29563
rect 36771 29529 36783 29563
rect 36725 29523 36783 29529
rect 28868 29464 34284 29492
rect 28868 29452 28874 29464
rect 34606 29452 34612 29504
rect 34664 29492 34670 29504
rect 35158 29492 35164 29504
rect 34664 29464 35164 29492
rect 34664 29452 34670 29464
rect 35158 29452 35164 29464
rect 35216 29452 35222 29504
rect 35250 29452 35256 29504
rect 35308 29492 35314 29504
rect 35529 29495 35587 29501
rect 35529 29492 35541 29495
rect 35308 29464 35541 29492
rect 35308 29452 35314 29464
rect 35529 29461 35541 29464
rect 35575 29492 35587 29495
rect 35618 29492 35624 29504
rect 35575 29464 35624 29492
rect 35575 29461 35587 29464
rect 35529 29455 35587 29461
rect 35618 29452 35624 29464
rect 35676 29452 35682 29504
rect 36740 29492 36768 29523
rect 36906 29520 36912 29572
rect 36964 29569 36970 29572
rect 36964 29563 36993 29569
rect 36981 29529 36993 29563
rect 36964 29523 36993 29529
rect 36964 29520 36970 29523
rect 37274 29492 37280 29504
rect 36740 29464 37280 29492
rect 37274 29452 37280 29464
rect 37332 29452 37338 29504
rect 37752 29492 37780 29591
rect 38654 29588 38660 29640
rect 38712 29628 38718 29640
rect 38841 29631 38899 29637
rect 38841 29628 38853 29631
rect 38712 29600 38853 29628
rect 38712 29588 38718 29600
rect 38841 29597 38853 29600
rect 38887 29597 38899 29631
rect 38841 29591 38899 29597
rect 38856 29560 38884 29591
rect 40126 29588 40132 29640
rect 40184 29628 40190 29640
rect 40313 29631 40371 29637
rect 40313 29628 40325 29631
rect 40184 29600 40325 29628
rect 40184 29588 40190 29600
rect 40313 29597 40325 29600
rect 40359 29628 40371 29631
rect 41064 29628 41276 29630
rect 41874 29628 41880 29640
rect 40359 29602 41880 29628
rect 40359 29600 41092 29602
rect 41248 29600 41880 29602
rect 40359 29597 40371 29600
rect 40313 29591 40371 29597
rect 41874 29588 41880 29600
rect 41932 29588 41938 29640
rect 43346 29588 43352 29640
rect 43404 29588 43410 29640
rect 43990 29628 43996 29640
rect 43951 29600 43996 29628
rect 43990 29588 43996 29600
rect 44048 29588 44054 29640
rect 44082 29588 44088 29640
rect 44140 29628 44146 29640
rect 44453 29631 44511 29637
rect 44453 29628 44465 29631
rect 44140 29600 44465 29628
rect 44140 29588 44146 29600
rect 44453 29597 44465 29600
rect 44499 29597 44511 29631
rect 45186 29628 45192 29640
rect 45147 29600 45192 29628
rect 44453 29591 44511 29597
rect 45186 29588 45192 29600
rect 45244 29588 45250 29640
rect 45278 29588 45284 29640
rect 45336 29628 45342 29640
rect 45480 29628 45508 29668
rect 46106 29656 46112 29708
rect 46164 29696 46170 29708
rect 46569 29699 46627 29705
rect 46569 29696 46581 29699
rect 46164 29668 46581 29696
rect 46164 29656 46170 29668
rect 46569 29665 46581 29668
rect 46615 29696 46627 29699
rect 46842 29696 46848 29708
rect 46615 29668 46848 29696
rect 46615 29665 46627 29668
rect 46569 29659 46627 29665
rect 46842 29656 46848 29668
rect 46900 29656 46906 29708
rect 47026 29696 47032 29708
rect 46987 29668 47032 29696
rect 47026 29656 47032 29668
rect 47084 29656 47090 29708
rect 47210 29656 47216 29708
rect 47268 29696 47274 29708
rect 50985 29699 51043 29705
rect 50985 29696 50997 29699
rect 47268 29668 50997 29696
rect 47268 29656 47274 29668
rect 50985 29665 50997 29668
rect 51031 29665 51043 29699
rect 51902 29696 51908 29708
rect 51863 29668 51908 29696
rect 50985 29659 51043 29665
rect 51902 29656 51908 29668
rect 51960 29656 51966 29708
rect 53558 29656 53564 29708
rect 53616 29696 53622 29708
rect 54128 29705 54156 29736
rect 56502 29724 56508 29736
rect 56560 29724 56566 29776
rect 56870 29724 56876 29776
rect 56928 29764 56934 29776
rect 56928 29736 57008 29764
rect 56928 29724 56934 29736
rect 54113 29699 54171 29705
rect 54113 29696 54125 29699
rect 53616 29668 54125 29696
rect 53616 29656 53622 29668
rect 54113 29665 54125 29668
rect 54159 29665 54171 29699
rect 54113 29659 54171 29665
rect 54481 29699 54539 29705
rect 54481 29665 54493 29699
rect 54527 29696 54539 29699
rect 54662 29696 54668 29708
rect 54527 29668 54668 29696
rect 54527 29665 54539 29668
rect 54481 29659 54539 29665
rect 54662 29656 54668 29668
rect 54720 29656 54726 29708
rect 55122 29656 55128 29708
rect 55180 29696 55186 29708
rect 56980 29705 57008 29736
rect 56965 29699 57023 29705
rect 55180 29668 56916 29696
rect 55180 29656 55186 29668
rect 45654 29631 45712 29637
rect 45654 29628 45666 29631
rect 45336 29600 45381 29628
rect 45480 29600 45666 29628
rect 45336 29588 45342 29600
rect 45654 29597 45666 29600
rect 45700 29597 45712 29631
rect 45654 29591 45712 29597
rect 46293 29631 46351 29637
rect 46293 29597 46305 29631
rect 46339 29628 46351 29631
rect 46658 29628 46664 29640
rect 46339 29600 46664 29628
rect 46339 29597 46351 29600
rect 46293 29591 46351 29597
rect 46658 29588 46664 29600
rect 46716 29588 46722 29640
rect 47305 29631 47363 29637
rect 47305 29597 47317 29631
rect 47351 29628 47363 29631
rect 47394 29628 47400 29640
rect 47351 29600 47400 29628
rect 47351 29597 47363 29600
rect 47305 29591 47363 29597
rect 47394 29588 47400 29600
rect 47452 29588 47458 29640
rect 47946 29588 47952 29640
rect 48004 29628 48010 29640
rect 48041 29631 48099 29637
rect 48041 29628 48053 29631
rect 48004 29600 48053 29628
rect 48004 29588 48010 29600
rect 48041 29597 48053 29600
rect 48087 29597 48099 29631
rect 48041 29591 48099 29597
rect 40037 29563 40095 29569
rect 40037 29560 40049 29563
rect 38856 29532 40049 29560
rect 40037 29529 40049 29532
rect 40083 29529 40095 29563
rect 40037 29523 40095 29529
rect 40221 29563 40279 29569
rect 40221 29529 40233 29563
rect 40267 29560 40279 29563
rect 41598 29560 41604 29572
rect 40267 29532 41604 29560
rect 40267 29529 40279 29532
rect 40221 29523 40279 29529
rect 41598 29520 41604 29532
rect 41656 29520 41662 29572
rect 41690 29520 41696 29572
rect 41748 29560 41754 29572
rect 42245 29563 42303 29569
rect 42245 29560 42257 29563
rect 41748 29532 42257 29560
rect 41748 29520 41754 29532
rect 42245 29529 42257 29532
rect 42291 29529 42303 29563
rect 42245 29523 42303 29529
rect 43806 29520 43812 29572
rect 43864 29560 43870 29572
rect 45462 29560 45468 29572
rect 43864 29532 45468 29560
rect 43864 29520 43870 29532
rect 45462 29520 45468 29532
rect 45520 29520 45526 29572
rect 45557 29563 45615 29569
rect 45557 29529 45569 29563
rect 45603 29560 45615 29563
rect 45738 29560 45744 29572
rect 45603 29532 45744 29560
rect 45603 29529 45615 29532
rect 45557 29523 45615 29529
rect 45738 29520 45744 29532
rect 45796 29520 45802 29572
rect 47854 29560 47860 29572
rect 47815 29532 47860 29560
rect 47854 29520 47860 29532
rect 47912 29520 47918 29572
rect 48056 29560 48084 29591
rect 48130 29588 48136 29640
rect 48188 29628 48194 29640
rect 48188 29600 48233 29628
rect 48188 29588 48194 29600
rect 48498 29588 48504 29640
rect 48556 29628 48562 29640
rect 48556 29600 49188 29628
rect 48556 29588 48562 29600
rect 48314 29560 48320 29572
rect 48056 29532 48320 29560
rect 48314 29520 48320 29532
rect 48372 29520 48378 29572
rect 49053 29563 49111 29569
rect 49053 29529 49065 29563
rect 49099 29529 49111 29563
rect 49160 29560 49188 29600
rect 50154 29588 50160 29640
rect 50212 29628 50218 29640
rect 50341 29631 50399 29637
rect 50341 29628 50353 29631
rect 50212 29600 50353 29628
rect 50212 29588 50218 29600
rect 50341 29597 50353 29600
rect 50387 29597 50399 29631
rect 50341 29591 50399 29597
rect 50525 29631 50583 29637
rect 50525 29597 50537 29631
rect 50571 29597 50583 29631
rect 50525 29591 50583 29597
rect 51997 29631 52055 29637
rect 51997 29597 52009 29631
rect 52043 29628 52055 29631
rect 52086 29628 52092 29640
rect 52043 29600 52092 29628
rect 52043 29597 52055 29600
rect 51997 29591 52055 29597
rect 49253 29563 49311 29569
rect 49253 29560 49265 29563
rect 49160 29532 49265 29560
rect 49053 29523 49111 29529
rect 49253 29529 49265 29532
rect 49299 29529 49311 29563
rect 49253 29523 49311 29529
rect 38930 29492 38936 29504
rect 37752 29464 38936 29492
rect 38930 29452 38936 29464
rect 38988 29452 38994 29504
rect 40313 29495 40371 29501
rect 40313 29461 40325 29495
rect 40359 29492 40371 29495
rect 40494 29492 40500 29504
rect 40359 29464 40500 29492
rect 40359 29461 40371 29464
rect 40313 29455 40371 29461
rect 40494 29452 40500 29464
rect 40552 29452 40558 29504
rect 41141 29495 41199 29501
rect 41141 29461 41153 29495
rect 41187 29492 41199 29495
rect 42518 29492 42524 29504
rect 41187 29464 42524 29492
rect 41187 29461 41199 29464
rect 41141 29455 41199 29461
rect 42518 29452 42524 29464
rect 42576 29492 42582 29504
rect 43070 29492 43076 29504
rect 42576 29464 43076 29492
rect 42576 29452 42582 29464
rect 43070 29452 43076 29464
rect 43128 29452 43134 29504
rect 47029 29495 47087 29501
rect 47029 29461 47041 29495
rect 47075 29492 47087 29495
rect 48682 29492 48688 29504
rect 47075 29464 48688 29492
rect 47075 29461 47087 29464
rect 47029 29455 47087 29461
rect 48682 29452 48688 29464
rect 48740 29452 48746 29504
rect 49068 29492 49096 29523
rect 49418 29520 49424 29572
rect 49476 29560 49482 29572
rect 50540 29560 50568 29591
rect 52086 29588 52092 29600
rect 52144 29588 52150 29640
rect 52822 29588 52828 29640
rect 52880 29588 52886 29640
rect 53098 29628 53104 29640
rect 53059 29600 53104 29628
rect 53098 29588 53104 29600
rect 53156 29588 53162 29640
rect 53193 29631 53251 29637
rect 53193 29597 53205 29631
rect 53239 29597 53251 29631
rect 53374 29628 53380 29640
rect 53335 29600 53380 29628
rect 53193 29591 53251 29597
rect 49476 29532 50568 29560
rect 52840 29560 52868 29588
rect 53208 29560 53236 29591
rect 53374 29588 53380 29600
rect 53432 29588 53438 29640
rect 53469 29631 53527 29637
rect 53469 29597 53481 29631
rect 53515 29628 53527 29631
rect 54205 29631 54263 29637
rect 53515 29600 53972 29628
rect 53515 29597 53527 29600
rect 53469 29591 53527 29597
rect 53558 29560 53564 29572
rect 52840 29532 53564 29560
rect 49476 29520 49482 29532
rect 53558 29520 53564 29532
rect 53616 29520 53622 29572
rect 49694 29492 49700 29504
rect 49068 29464 49700 29492
rect 49694 29452 49700 29464
rect 49752 29452 49758 29504
rect 49786 29452 49792 29504
rect 49844 29492 49850 29504
rect 50433 29495 50491 29501
rect 50433 29492 50445 29495
rect 49844 29464 50445 29492
rect 49844 29452 49850 29464
rect 50433 29461 50445 29464
rect 50479 29461 50491 29495
rect 50433 29455 50491 29461
rect 52365 29495 52423 29501
rect 52365 29461 52377 29495
rect 52411 29492 52423 29495
rect 52822 29492 52828 29504
rect 52411 29464 52828 29492
rect 52411 29461 52423 29464
rect 52365 29455 52423 29461
rect 52822 29452 52828 29464
rect 52880 29452 52886 29504
rect 52917 29495 52975 29501
rect 52917 29461 52929 29495
rect 52963 29492 52975 29495
rect 53282 29492 53288 29504
rect 52963 29464 53288 29492
rect 52963 29461 52975 29464
rect 52917 29455 52975 29461
rect 53282 29452 53288 29464
rect 53340 29452 53346 29504
rect 53944 29501 53972 29600
rect 54205 29597 54217 29631
rect 54251 29628 54263 29631
rect 55490 29628 55496 29640
rect 54251 29600 55496 29628
rect 54251 29597 54263 29600
rect 54205 29591 54263 29597
rect 55490 29588 55496 29600
rect 55548 29588 55554 29640
rect 55582 29588 55588 29640
rect 55640 29628 55646 29640
rect 55677 29631 55735 29637
rect 55677 29628 55689 29631
rect 55640 29600 55689 29628
rect 55640 29588 55646 29600
rect 55677 29597 55689 29600
rect 55723 29597 55735 29631
rect 55677 29591 55735 29597
rect 55766 29588 55772 29640
rect 55824 29628 55830 29640
rect 56042 29628 56048 29640
rect 55824 29600 55869 29628
rect 56003 29600 56048 29628
rect 55824 29588 55830 29600
rect 56042 29588 56048 29600
rect 56100 29588 56106 29640
rect 56888 29637 56916 29668
rect 56965 29665 56977 29699
rect 57011 29665 57023 29699
rect 57238 29696 57244 29708
rect 57199 29668 57244 29696
rect 56965 29659 57023 29665
rect 57238 29656 57244 29668
rect 57296 29656 57302 29708
rect 56873 29631 56931 29637
rect 56873 29597 56885 29631
rect 56919 29597 56931 29631
rect 56873 29591 56931 29597
rect 57974 29588 57980 29640
rect 58032 29628 58038 29640
rect 58069 29631 58127 29637
rect 58069 29628 58081 29631
rect 58032 29600 58081 29628
rect 58032 29588 58038 29600
rect 58069 29597 58081 29600
rect 58115 29597 58127 29631
rect 58069 29591 58127 29597
rect 54573 29563 54631 29569
rect 54573 29529 54585 29563
rect 54619 29560 54631 29563
rect 55306 29560 55312 29572
rect 54619 29532 55312 29560
rect 54619 29529 54631 29532
rect 54573 29523 54631 29529
rect 55306 29520 55312 29532
rect 55364 29560 55370 29572
rect 56137 29563 56195 29569
rect 56137 29560 56149 29563
rect 55364 29532 56149 29560
rect 55364 29520 55370 29532
rect 56137 29529 56149 29532
rect 56183 29560 56195 29563
rect 56410 29560 56416 29572
rect 56183 29532 56416 29560
rect 56183 29529 56195 29532
rect 56137 29523 56195 29529
rect 56410 29520 56416 29532
rect 56468 29520 56474 29572
rect 53929 29495 53987 29501
rect 53929 29461 53941 29495
rect 53975 29461 53987 29495
rect 55490 29492 55496 29504
rect 55451 29464 55496 29492
rect 53929 29455 53987 29461
rect 55490 29452 55496 29464
rect 55548 29452 55554 29504
rect 58250 29492 58256 29504
rect 58211 29464 58256 29492
rect 58250 29452 58256 29464
rect 58308 29452 58314 29504
rect 1104 29402 58880 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 58880 29402
rect 1104 29328 58880 29350
rect 30190 29288 30196 29300
rect 30151 29260 30196 29288
rect 30190 29248 30196 29260
rect 30248 29248 30254 29300
rect 32677 29291 32735 29297
rect 32677 29257 32689 29291
rect 32723 29288 32735 29291
rect 32766 29288 32772 29300
rect 32723 29260 32772 29288
rect 32723 29257 32735 29260
rect 32677 29251 32735 29257
rect 32766 29248 32772 29260
rect 32824 29248 32830 29300
rect 36814 29288 36820 29300
rect 36096 29260 36820 29288
rect 30101 29155 30159 29161
rect 30101 29121 30113 29155
rect 30147 29152 30159 29155
rect 30837 29155 30895 29161
rect 30837 29152 30849 29155
rect 30147 29124 30849 29152
rect 30147 29121 30159 29124
rect 30101 29115 30159 29121
rect 30837 29121 30849 29124
rect 30883 29152 30895 29155
rect 31754 29152 31760 29164
rect 30883 29124 31760 29152
rect 30883 29121 30895 29124
rect 30837 29115 30895 29121
rect 31754 29112 31760 29124
rect 31812 29152 31818 29164
rect 32585 29155 32643 29161
rect 31812 29124 31857 29152
rect 31812 29112 31818 29124
rect 32585 29121 32597 29155
rect 32631 29152 32643 29155
rect 32858 29152 32864 29164
rect 32631 29124 32864 29152
rect 32631 29121 32643 29124
rect 32585 29115 32643 29121
rect 32858 29112 32864 29124
rect 32916 29112 32922 29164
rect 33410 29152 33416 29164
rect 33371 29124 33416 29152
rect 33410 29112 33416 29124
rect 33468 29112 33474 29164
rect 34790 29112 34796 29164
rect 34848 29112 34854 29164
rect 36096 29161 36124 29260
rect 36814 29248 36820 29260
rect 36872 29248 36878 29300
rect 36909 29291 36967 29297
rect 36909 29257 36921 29291
rect 36955 29288 36967 29291
rect 37366 29288 37372 29300
rect 36955 29260 37372 29288
rect 36955 29257 36967 29260
rect 36909 29251 36967 29257
rect 37366 29248 37372 29260
rect 37424 29248 37430 29300
rect 37642 29248 37648 29300
rect 37700 29288 37706 29300
rect 37829 29291 37887 29297
rect 37829 29288 37841 29291
rect 37700 29260 37841 29288
rect 37700 29248 37706 29260
rect 37829 29257 37841 29260
rect 37875 29257 37887 29291
rect 39206 29288 39212 29300
rect 39167 29260 39212 29288
rect 37829 29251 37887 29257
rect 39206 29248 39212 29260
rect 39264 29248 39270 29300
rect 39853 29291 39911 29297
rect 39853 29288 39865 29291
rect 39316 29260 39865 29288
rect 36354 29180 36360 29232
rect 36412 29220 36418 29232
rect 39316 29220 39344 29260
rect 39853 29257 39865 29260
rect 39899 29257 39911 29291
rect 39853 29251 39911 29257
rect 40034 29248 40040 29300
rect 40092 29288 40098 29300
rect 40092 29260 40172 29288
rect 40092 29248 40098 29260
rect 40144 29229 40172 29260
rect 41138 29248 41144 29300
rect 41196 29288 41202 29300
rect 41690 29288 41696 29300
rect 41196 29260 41552 29288
rect 41651 29260 41696 29288
rect 41196 29248 41202 29260
rect 36412 29192 39344 29220
rect 40129 29223 40187 29229
rect 36412 29180 36418 29192
rect 40129 29189 40141 29223
rect 40175 29189 40187 29223
rect 40129 29183 40187 29189
rect 40221 29223 40279 29229
rect 40221 29189 40233 29223
rect 40267 29220 40279 29223
rect 40770 29220 40776 29232
rect 40267 29192 40776 29220
rect 40267 29189 40279 29192
rect 40221 29183 40279 29189
rect 40770 29180 40776 29192
rect 40828 29180 40834 29232
rect 40862 29180 40868 29232
rect 40920 29220 40926 29232
rect 41414 29220 41420 29232
rect 40920 29192 41420 29220
rect 40920 29180 40926 29192
rect 41414 29180 41420 29192
rect 41472 29180 41478 29232
rect 36000 29155 36058 29161
rect 35898 29145 35956 29151
rect 35898 29111 35910 29145
rect 35944 29111 35956 29145
rect 36000 29121 36012 29155
rect 36046 29121 36058 29155
rect 36000 29115 36058 29121
rect 36094 29155 36152 29161
rect 36094 29121 36106 29155
rect 36140 29121 36152 29155
rect 36094 29115 36152 29121
rect 36219 29155 36277 29161
rect 36219 29121 36231 29155
rect 36265 29152 36277 29155
rect 36906 29152 36912 29164
rect 36265 29124 36912 29152
rect 36265 29121 36277 29124
rect 36219 29115 36277 29121
rect 35898 29105 35956 29111
rect 33686 29084 33692 29096
rect 33647 29056 33692 29084
rect 33686 29044 33692 29056
rect 33744 29044 33750 29096
rect 33778 29044 33784 29096
rect 33836 29084 33842 29096
rect 35713 29087 35771 29093
rect 35713 29084 35725 29087
rect 33836 29056 35725 29084
rect 33836 29044 33842 29056
rect 35713 29053 35725 29056
rect 35759 29053 35771 29087
rect 35713 29047 35771 29053
rect 35912 29028 35940 29105
rect 36005 29028 36033 29115
rect 36906 29112 36912 29124
rect 36964 29112 36970 29164
rect 37550 29112 37556 29164
rect 37608 29152 37614 29164
rect 38381 29155 38439 29161
rect 38381 29152 38393 29155
rect 37608 29124 38393 29152
rect 37608 29112 37614 29124
rect 38381 29121 38393 29124
rect 38427 29121 38439 29155
rect 38838 29152 38844 29164
rect 38799 29124 38844 29152
rect 38381 29115 38439 29121
rect 38838 29112 38844 29124
rect 38896 29112 38902 29164
rect 39025 29155 39083 29161
rect 39025 29121 39037 29155
rect 39071 29121 39083 29155
rect 39025 29115 39083 29121
rect 36354 29084 36360 29096
rect 36315 29056 36360 29084
rect 36354 29044 36360 29056
rect 36412 29044 36418 29096
rect 38105 29087 38163 29093
rect 38105 29053 38117 29087
rect 38151 29084 38163 29087
rect 38562 29084 38568 29096
rect 38151 29056 38568 29084
rect 38151 29053 38163 29056
rect 38105 29047 38163 29053
rect 38562 29044 38568 29056
rect 38620 29044 38626 29096
rect 38930 29044 38936 29096
rect 38988 29084 38994 29096
rect 39040 29084 39068 29115
rect 39942 29112 39948 29164
rect 40000 29152 40006 29164
rect 40037 29155 40095 29161
rect 40037 29152 40049 29155
rect 40000 29124 40049 29152
rect 40000 29112 40006 29124
rect 40037 29121 40049 29124
rect 40083 29121 40095 29155
rect 40037 29115 40095 29121
rect 40310 29112 40316 29164
rect 40368 29161 40374 29164
rect 40368 29155 40417 29161
rect 40368 29121 40371 29155
rect 40405 29121 40417 29155
rect 40368 29115 40417 29121
rect 40368 29112 40374 29115
rect 40494 29112 40500 29164
rect 40552 29152 40558 29164
rect 41046 29152 41052 29164
rect 40552 29124 40597 29152
rect 41007 29124 41052 29152
rect 40552 29112 40558 29124
rect 41046 29112 41052 29124
rect 41104 29112 41110 29164
rect 41230 29161 41236 29164
rect 41207 29155 41236 29161
rect 41207 29121 41219 29155
rect 41207 29115 41236 29121
rect 41230 29112 41236 29115
rect 41288 29112 41294 29164
rect 41524 29161 41552 29260
rect 41690 29248 41696 29260
rect 41748 29248 41754 29300
rect 43346 29248 43352 29300
rect 43404 29288 43410 29300
rect 43441 29291 43499 29297
rect 43441 29288 43453 29291
rect 43404 29260 43453 29288
rect 43404 29248 43410 29260
rect 43441 29257 43453 29260
rect 43487 29257 43499 29291
rect 49878 29288 49884 29300
rect 43441 29251 43499 29257
rect 46768 29260 49884 29288
rect 41874 29180 41880 29232
rect 41932 29220 41938 29232
rect 44082 29220 44088 29232
rect 41932 29192 42932 29220
rect 41932 29180 41938 29192
rect 42904 29161 42932 29192
rect 43548 29192 44088 29220
rect 41325 29155 41383 29161
rect 41325 29121 41337 29155
rect 41371 29121 41383 29155
rect 41325 29115 41383 29121
rect 41509 29155 41567 29161
rect 41509 29121 41521 29155
rect 41555 29121 41567 29155
rect 41509 29115 41567 29121
rect 42613 29155 42671 29161
rect 42613 29121 42625 29155
rect 42659 29121 42671 29155
rect 42613 29115 42671 29121
rect 42797 29155 42855 29161
rect 42797 29121 42809 29155
rect 42843 29121 42855 29155
rect 42797 29115 42855 29121
rect 42889 29155 42947 29161
rect 42889 29121 42901 29155
rect 42935 29121 42947 29155
rect 42889 29115 42947 29121
rect 38988 29056 40172 29084
rect 38988 29044 38994 29056
rect 35158 29016 35164 29028
rect 35119 28988 35164 29016
rect 35158 28976 35164 28988
rect 35216 29016 35222 29028
rect 35802 29016 35808 29028
rect 35216 28988 35808 29016
rect 35216 28976 35222 28988
rect 35802 28976 35808 28988
rect 35860 28976 35866 29028
rect 35894 28976 35900 29028
rect 35952 28976 35958 29028
rect 35986 28976 35992 29028
rect 36044 29016 36050 29028
rect 39114 29016 39120 29028
rect 36044 28988 39120 29016
rect 36044 28976 36050 28988
rect 39114 28976 39120 28988
rect 39172 28976 39178 29028
rect 40144 28994 40172 29056
rect 40770 29044 40776 29096
rect 40828 29084 40834 29096
rect 41340 29084 41368 29115
rect 42628 29084 42656 29115
rect 40828 29056 41368 29084
rect 41432 29056 42656 29084
rect 40828 29044 40834 29056
rect 40144 28966 40382 28994
rect 31662 28948 31668 28960
rect 31623 28920 31668 28948
rect 31662 28908 31668 28920
rect 31720 28908 31726 28960
rect 35250 28908 35256 28960
rect 35308 28948 35314 28960
rect 35710 28948 35716 28960
rect 35308 28920 35716 28948
rect 35308 28908 35314 28920
rect 35710 28908 35716 28920
rect 35768 28908 35774 28960
rect 36078 28908 36084 28960
rect 36136 28948 36142 28960
rect 37826 28948 37832 28960
rect 36136 28920 37832 28948
rect 36136 28908 36142 28920
rect 37826 28908 37832 28920
rect 37884 28908 37890 28960
rect 38289 28951 38347 28957
rect 38289 28917 38301 28951
rect 38335 28948 38347 28951
rect 40034 28948 40040 28960
rect 38335 28920 40040 28948
rect 38335 28917 38347 28920
rect 38289 28911 38347 28917
rect 40034 28908 40040 28920
rect 40092 28908 40098 28960
rect 40354 28948 40382 28966
rect 41432 28948 41460 29056
rect 42812 29016 42840 29115
rect 42978 29112 42984 29164
rect 43036 29152 43042 29164
rect 43548 29161 43576 29192
rect 44082 29180 44088 29192
rect 44140 29180 44146 29232
rect 46198 29180 46204 29232
rect 46256 29220 46262 29232
rect 46768 29220 46796 29260
rect 49878 29248 49884 29260
rect 49936 29248 49942 29300
rect 55214 29288 55220 29300
rect 53852 29260 55220 29288
rect 46256 29192 46796 29220
rect 46256 29180 46262 29192
rect 43533 29155 43591 29161
rect 43533 29152 43545 29155
rect 43036 29124 43545 29152
rect 43036 29112 43042 29124
rect 43533 29121 43545 29124
rect 43579 29121 43591 29155
rect 43533 29115 43591 29121
rect 43898 29112 43904 29164
rect 43956 29152 43962 29164
rect 43956 29124 44404 29152
rect 43956 29112 43962 29124
rect 43806 29044 43812 29096
rect 43864 29084 43870 29096
rect 44085 29087 44143 29093
rect 44085 29084 44097 29087
rect 43864 29056 44097 29084
rect 43864 29044 43870 29056
rect 44085 29053 44097 29056
rect 44131 29053 44143 29087
rect 44266 29084 44272 29096
rect 44227 29056 44272 29084
rect 44085 29047 44143 29053
rect 44266 29044 44272 29056
rect 44324 29044 44330 29096
rect 44376 29084 44404 29124
rect 45094 29112 45100 29164
rect 45152 29161 45158 29164
rect 45152 29155 45180 29161
rect 45168 29121 45180 29155
rect 46106 29152 46112 29164
rect 45152 29115 45180 29121
rect 45848 29124 46112 29152
rect 45152 29112 45158 29115
rect 45005 29087 45063 29093
rect 45005 29084 45017 29087
rect 44376 29056 45017 29084
rect 45005 29053 45017 29056
rect 45051 29053 45063 29087
rect 45005 29047 45063 29053
rect 45281 29087 45339 29093
rect 45281 29053 45293 29087
rect 45327 29084 45339 29087
rect 45848 29084 45876 29124
rect 46106 29112 46112 29124
rect 46164 29112 46170 29164
rect 46290 29112 46296 29164
rect 46348 29152 46354 29164
rect 46768 29161 46796 29192
rect 47670 29180 47676 29232
rect 47728 29220 47734 29232
rect 48133 29223 48191 29229
rect 48133 29220 48145 29223
rect 47728 29192 48145 29220
rect 47728 29180 47734 29192
rect 48133 29189 48145 29192
rect 48179 29189 48191 29223
rect 50154 29220 50160 29232
rect 48133 29183 48191 29189
rect 49436 29192 50160 29220
rect 46661 29155 46719 29161
rect 46661 29152 46673 29155
rect 46348 29124 46673 29152
rect 46348 29112 46354 29124
rect 46661 29121 46673 29124
rect 46707 29121 46719 29155
rect 46661 29115 46719 29121
rect 46753 29155 46811 29161
rect 46753 29121 46765 29155
rect 46799 29121 46811 29155
rect 46934 29152 46940 29164
rect 46895 29124 46940 29152
rect 46753 29115 46811 29121
rect 46934 29112 46940 29124
rect 46992 29112 46998 29164
rect 47029 29155 47087 29161
rect 47029 29121 47041 29155
rect 47075 29152 47087 29155
rect 47486 29152 47492 29164
rect 47075 29124 47492 29152
rect 47075 29121 47087 29124
rect 47029 29115 47087 29121
rect 47486 29112 47492 29124
rect 47544 29112 47550 29164
rect 47946 29161 47952 29164
rect 47772 29155 47830 29161
rect 47772 29121 47784 29155
rect 47818 29121 47830 29155
rect 47772 29115 47830 29121
rect 47913 29155 47952 29161
rect 47913 29121 47925 29155
rect 47913 29115 47952 29121
rect 45327 29056 45876 29084
rect 45925 29087 45983 29093
rect 45327 29053 45339 29056
rect 45281 29047 45339 29053
rect 45925 29053 45937 29087
rect 45971 29084 45983 29087
rect 46474 29084 46480 29096
rect 45971 29056 46480 29084
rect 45971 29053 45983 29056
rect 45925 29047 45983 29053
rect 46474 29044 46480 29056
rect 46532 29044 46538 29096
rect 46842 29044 46848 29096
rect 46900 29084 46906 29096
rect 47780 29084 47808 29115
rect 47946 29112 47952 29115
rect 48004 29112 48010 29164
rect 48314 29161 48320 29164
rect 48041 29155 48099 29161
rect 48041 29121 48053 29155
rect 48087 29121 48099 29155
rect 48041 29115 48099 29121
rect 48271 29155 48320 29161
rect 48271 29121 48283 29155
rect 48317 29121 48320 29155
rect 48271 29115 48320 29121
rect 48056 29084 48084 29115
rect 48314 29112 48320 29115
rect 48372 29112 48378 29164
rect 49436 29161 49464 29192
rect 50154 29180 50160 29192
rect 50212 29180 50218 29232
rect 53852 29229 53880 29260
rect 55214 29248 55220 29260
rect 55272 29248 55278 29300
rect 58161 29291 58219 29297
rect 58161 29257 58173 29291
rect 58207 29288 58219 29291
rect 58342 29288 58348 29300
rect 58207 29260 58348 29288
rect 58207 29257 58219 29260
rect 58161 29251 58219 29257
rect 58342 29248 58348 29260
rect 58400 29248 58406 29300
rect 53837 29223 53895 29229
rect 53837 29189 53849 29223
rect 53883 29189 53895 29223
rect 53837 29183 53895 29189
rect 54662 29180 54668 29232
rect 54720 29220 54726 29232
rect 55582 29220 55588 29232
rect 54720 29192 55588 29220
rect 54720 29180 54726 29192
rect 49421 29155 49479 29161
rect 49421 29121 49433 29155
rect 49467 29121 49479 29155
rect 49421 29115 49479 29121
rect 49510 29112 49516 29164
rect 49568 29152 49574 29164
rect 49694 29152 49700 29164
rect 49568 29124 49613 29152
rect 49655 29124 49700 29152
rect 49568 29112 49574 29124
rect 49694 29112 49700 29124
rect 49752 29112 49758 29164
rect 49789 29155 49847 29161
rect 49789 29121 49801 29155
rect 49835 29152 49847 29155
rect 49878 29152 49884 29164
rect 49835 29124 49884 29152
rect 49835 29121 49847 29124
rect 49789 29115 49847 29121
rect 49878 29112 49884 29124
rect 49936 29112 49942 29164
rect 50614 29112 50620 29164
rect 50672 29152 50678 29164
rect 50709 29155 50767 29161
rect 50709 29152 50721 29155
rect 50672 29124 50721 29152
rect 50672 29112 50678 29124
rect 50709 29121 50721 29124
rect 50755 29121 50767 29155
rect 51350 29152 51356 29164
rect 50709 29115 50767 29121
rect 50816 29124 51356 29152
rect 50816 29093 50844 29124
rect 51350 29112 51356 29124
rect 51408 29112 51414 29164
rect 51718 29112 51724 29164
rect 51776 29152 51782 29164
rect 51905 29155 51963 29161
rect 51905 29152 51917 29155
rect 51776 29124 51917 29152
rect 51776 29112 51782 29124
rect 51905 29121 51917 29124
rect 51951 29121 51963 29155
rect 51905 29115 51963 29121
rect 52822 29112 52828 29164
rect 52880 29152 52886 29164
rect 53009 29155 53067 29161
rect 53009 29152 53021 29155
rect 52880 29124 53021 29152
rect 52880 29112 52886 29124
rect 53009 29121 53021 29124
rect 53055 29121 53067 29155
rect 53009 29115 53067 29121
rect 53193 29155 53251 29161
rect 53193 29121 53205 29155
rect 53239 29152 53251 29155
rect 53466 29152 53472 29164
rect 53239 29124 53472 29152
rect 53239 29121 53251 29124
rect 53193 29115 53251 29121
rect 53466 29112 53472 29124
rect 53524 29112 53530 29164
rect 54021 29155 54079 29161
rect 54021 29121 54033 29155
rect 54067 29152 54079 29155
rect 54386 29152 54392 29164
rect 54067 29124 54392 29152
rect 54067 29121 54079 29124
rect 54021 29115 54079 29121
rect 54386 29112 54392 29124
rect 54444 29112 54450 29164
rect 55232 29161 55260 29192
rect 55582 29180 55588 29192
rect 55640 29180 55646 29232
rect 56686 29180 56692 29232
rect 56744 29220 56750 29232
rect 56965 29223 57023 29229
rect 56965 29220 56977 29223
rect 56744 29192 56977 29220
rect 56744 29180 56750 29192
rect 56965 29189 56977 29192
rect 57011 29189 57023 29223
rect 56965 29183 57023 29189
rect 55125 29155 55183 29161
rect 55125 29152 55137 29155
rect 54496 29124 55137 29152
rect 46900 29056 47808 29084
rect 47872 29056 48084 29084
rect 50801 29087 50859 29093
rect 46900 29044 46906 29056
rect 47872 29028 47900 29056
rect 50801 29053 50813 29087
rect 50847 29053 50859 29087
rect 50801 29047 50859 29053
rect 51077 29087 51135 29093
rect 51077 29053 51089 29087
rect 51123 29084 51135 29087
rect 51813 29087 51871 29093
rect 51813 29084 51825 29087
rect 51123 29056 51825 29084
rect 51123 29053 51135 29056
rect 51077 29047 51135 29053
rect 51813 29053 51825 29056
rect 51859 29053 51871 29087
rect 51813 29047 51871 29053
rect 53098 29044 53104 29096
rect 53156 29084 53162 29096
rect 54496 29084 54524 29124
rect 55125 29121 55137 29124
rect 55171 29121 55183 29155
rect 55125 29115 55183 29121
rect 55217 29155 55275 29161
rect 55217 29121 55229 29155
rect 55263 29121 55275 29155
rect 55398 29152 55404 29164
rect 55359 29124 55404 29152
rect 55217 29115 55275 29121
rect 53156 29056 54524 29084
rect 55140 29084 55168 29115
rect 55398 29112 55404 29124
rect 55456 29112 55462 29164
rect 55490 29112 55496 29164
rect 55548 29152 55554 29164
rect 55950 29152 55956 29164
rect 55548 29124 55593 29152
rect 55911 29124 55956 29152
rect 55548 29112 55554 29124
rect 55950 29112 55956 29124
rect 56008 29112 56014 29164
rect 56045 29155 56103 29161
rect 56045 29121 56057 29155
rect 56091 29121 56103 29155
rect 56045 29115 56103 29121
rect 55416 29084 55444 29112
rect 56060 29084 56088 29115
rect 56134 29112 56140 29164
rect 56192 29152 56198 29164
rect 56229 29155 56287 29161
rect 56229 29152 56241 29155
rect 56192 29124 56241 29152
rect 56192 29112 56198 29124
rect 56229 29121 56241 29124
rect 56275 29121 56287 29155
rect 56229 29115 56287 29121
rect 56321 29155 56379 29161
rect 56321 29121 56333 29155
rect 56367 29121 56379 29155
rect 57330 29152 57336 29164
rect 57291 29124 57336 29152
rect 56321 29115 56379 29121
rect 55140 29056 55214 29084
rect 55416 29056 56088 29084
rect 53156 29044 53162 29056
rect 44726 29016 44732 29028
rect 41800 28988 42840 29016
rect 44687 28988 44732 29016
rect 40354 28920 41460 28948
rect 41598 28908 41604 28960
rect 41656 28948 41662 28960
rect 41800 28948 41828 28988
rect 44726 28976 44732 28988
rect 44784 28976 44790 29028
rect 47854 28976 47860 29028
rect 47912 29016 47918 29028
rect 48130 29016 48136 29028
rect 47912 28988 48136 29016
rect 47912 28976 47918 28988
rect 48130 28976 48136 28988
rect 48188 28976 48194 29028
rect 55186 29016 55214 29056
rect 56336 29016 56364 29115
rect 57330 29112 57336 29124
rect 57388 29112 57394 29164
rect 55186 28988 56364 29016
rect 42702 28948 42708 28960
rect 41656 28920 41828 28948
rect 42663 28920 42708 28948
rect 41656 28908 41662 28920
rect 42702 28908 42708 28920
rect 42760 28908 42766 28960
rect 46477 28951 46535 28957
rect 46477 28917 46489 28951
rect 46523 28948 46535 28951
rect 47026 28948 47032 28960
rect 46523 28920 47032 28948
rect 46523 28917 46535 28920
rect 46477 28911 46535 28917
rect 47026 28908 47032 28920
rect 47084 28908 47090 28960
rect 48409 28951 48467 28957
rect 48409 28917 48421 28951
rect 48455 28948 48467 28951
rect 48774 28948 48780 28960
rect 48455 28920 48780 28948
rect 48455 28917 48467 28920
rect 48409 28911 48467 28917
rect 48774 28908 48780 28920
rect 48832 28908 48838 28960
rect 49142 28908 49148 28960
rect 49200 28948 49206 28960
rect 49237 28951 49295 28957
rect 49237 28948 49249 28951
rect 49200 28920 49249 28948
rect 49200 28908 49206 28920
rect 49237 28917 49249 28920
rect 49283 28917 49295 28951
rect 49237 28911 49295 28917
rect 49326 28908 49332 28960
rect 49384 28948 49390 28960
rect 50798 28948 50804 28960
rect 49384 28920 50804 28948
rect 49384 28908 49390 28920
rect 50798 28908 50804 28920
rect 50856 28908 50862 28960
rect 51534 28948 51540 28960
rect 51495 28920 51540 28948
rect 51534 28908 51540 28920
rect 51592 28908 51598 28960
rect 53101 28951 53159 28957
rect 53101 28917 53113 28951
rect 53147 28948 53159 28951
rect 53466 28948 53472 28960
rect 53147 28920 53472 28948
rect 53147 28917 53159 28920
rect 53101 28911 53159 28917
rect 53466 28908 53472 28920
rect 53524 28908 53530 28960
rect 53650 28948 53656 28960
rect 53611 28920 53656 28948
rect 53650 28908 53656 28920
rect 53708 28908 53714 28960
rect 54846 28908 54852 28960
rect 54904 28948 54910 28960
rect 54941 28951 54999 28957
rect 54941 28948 54953 28951
rect 54904 28920 54953 28948
rect 54904 28908 54910 28920
rect 54941 28917 54953 28920
rect 54987 28917 54999 28951
rect 54941 28911 54999 28917
rect 55582 28908 55588 28960
rect 55640 28948 55646 28960
rect 56505 28951 56563 28957
rect 56505 28948 56517 28951
rect 55640 28920 56517 28948
rect 55640 28908 55646 28920
rect 56505 28917 56517 28920
rect 56551 28917 56563 28951
rect 56505 28911 56563 28917
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 30837 28747 30895 28753
rect 30837 28713 30849 28747
rect 30883 28744 30895 28747
rect 31202 28744 31208 28756
rect 30883 28716 31208 28744
rect 30883 28713 30895 28716
rect 30837 28707 30895 28713
rect 31202 28704 31208 28716
rect 31260 28744 31266 28756
rect 34330 28744 34336 28756
rect 31260 28716 34100 28744
rect 34291 28716 34336 28744
rect 31260 28704 31266 28716
rect 34072 28676 34100 28716
rect 34330 28704 34336 28716
rect 34388 28744 34394 28756
rect 34606 28744 34612 28756
rect 34388 28716 34612 28744
rect 34388 28704 34394 28716
rect 34606 28704 34612 28716
rect 34664 28704 34670 28756
rect 34790 28704 34796 28756
rect 34848 28744 34854 28756
rect 34977 28747 35035 28753
rect 34977 28744 34989 28747
rect 34848 28716 34989 28744
rect 34848 28704 34854 28716
rect 34977 28713 34989 28716
rect 35023 28713 35035 28747
rect 34977 28707 35035 28713
rect 36817 28747 36875 28753
rect 36817 28713 36829 28747
rect 36863 28744 36875 28747
rect 36906 28744 36912 28756
rect 36863 28716 36912 28744
rect 36863 28713 36875 28716
rect 36817 28707 36875 28713
rect 36906 28704 36912 28716
rect 36964 28704 36970 28756
rect 37185 28747 37243 28753
rect 37185 28713 37197 28747
rect 37231 28744 37243 28747
rect 37274 28744 37280 28756
rect 37231 28716 37280 28744
rect 37231 28713 37243 28716
rect 37185 28707 37243 28713
rect 37274 28704 37280 28716
rect 37332 28704 37338 28756
rect 40034 28744 40040 28756
rect 39995 28716 40040 28744
rect 40034 28704 40040 28716
rect 40092 28704 40098 28756
rect 40218 28704 40224 28756
rect 40276 28744 40282 28756
rect 40405 28747 40463 28753
rect 40405 28744 40417 28747
rect 40276 28716 40417 28744
rect 40276 28704 40282 28716
rect 40405 28713 40417 28716
rect 40451 28713 40463 28747
rect 45186 28744 45192 28756
rect 40405 28707 40463 28713
rect 41340 28716 43392 28744
rect 45147 28716 45192 28744
rect 36354 28676 36360 28688
rect 34072 28648 36360 28676
rect 36354 28636 36360 28648
rect 36412 28636 36418 28688
rect 38562 28676 38568 28688
rect 37108 28648 38568 28676
rect 32306 28568 32312 28620
rect 32364 28608 32370 28620
rect 32585 28611 32643 28617
rect 32585 28608 32597 28611
rect 32364 28580 32597 28608
rect 32364 28568 32370 28580
rect 32585 28577 32597 28580
rect 32631 28577 32643 28611
rect 32585 28571 32643 28577
rect 33686 28568 33692 28620
rect 33744 28608 33750 28620
rect 35713 28611 35771 28617
rect 35713 28608 35725 28611
rect 33744 28580 35725 28608
rect 33744 28568 33750 28580
rect 35713 28577 35725 28580
rect 35759 28577 35771 28611
rect 35713 28571 35771 28577
rect 35802 28568 35808 28620
rect 35860 28608 35866 28620
rect 37108 28617 37136 28648
rect 38562 28636 38568 28648
rect 38620 28636 38626 28688
rect 39666 28636 39672 28688
rect 39724 28676 39730 28688
rect 41340 28676 41368 28716
rect 39724 28648 41368 28676
rect 41432 28648 42840 28676
rect 39724 28636 39730 28648
rect 37093 28611 37151 28617
rect 35860 28580 36400 28608
rect 35860 28568 35866 28580
rect 32858 28500 32864 28552
rect 32916 28540 32922 28552
rect 33045 28543 33103 28549
rect 33045 28540 33057 28543
rect 32916 28512 33057 28540
rect 32916 28500 32922 28512
rect 33045 28509 33057 28512
rect 33091 28509 33103 28543
rect 33045 28503 33103 28509
rect 34790 28500 34796 28552
rect 34848 28540 34854 28552
rect 35069 28543 35127 28549
rect 35069 28540 35081 28543
rect 34848 28512 35081 28540
rect 34848 28500 34854 28512
rect 35069 28509 35081 28512
rect 35115 28540 35127 28543
rect 35434 28540 35440 28552
rect 35115 28512 35440 28540
rect 35115 28509 35127 28512
rect 35069 28503 35127 28509
rect 35434 28500 35440 28512
rect 35492 28500 35498 28552
rect 35894 28540 35900 28552
rect 35807 28512 35900 28540
rect 35894 28500 35900 28512
rect 35952 28500 35958 28552
rect 35986 28500 35992 28552
rect 36044 28540 36050 28552
rect 36372 28549 36400 28580
rect 37093 28577 37105 28611
rect 37139 28577 37151 28611
rect 37093 28571 37151 28577
rect 37182 28568 37188 28620
rect 37240 28608 37246 28620
rect 38013 28611 38071 28617
rect 38013 28608 38025 28611
rect 37240 28580 38025 28608
rect 37240 28568 37246 28580
rect 38013 28577 38025 28580
rect 38059 28577 38071 28611
rect 38013 28571 38071 28577
rect 38378 28568 38384 28620
rect 38436 28608 38442 28620
rect 41432 28608 41460 28648
rect 42702 28608 42708 28620
rect 38436 28580 41460 28608
rect 41524 28580 42708 28608
rect 38436 28568 38442 28580
rect 36357 28543 36415 28549
rect 36044 28512 36089 28540
rect 36044 28500 36050 28512
rect 36357 28509 36369 28543
rect 36403 28509 36415 28543
rect 36357 28503 36415 28509
rect 37369 28543 37427 28549
rect 37369 28509 37381 28543
rect 37415 28540 37427 28543
rect 37550 28540 37556 28552
rect 37415 28512 37556 28540
rect 37415 28509 37427 28512
rect 37369 28503 37427 28509
rect 37550 28500 37556 28512
rect 37608 28500 37614 28552
rect 38102 28540 38108 28552
rect 38063 28512 38108 28540
rect 38102 28500 38108 28512
rect 38160 28500 38166 28552
rect 38194 28500 38200 28552
rect 38252 28540 38258 28552
rect 38252 28512 38297 28540
rect 38252 28500 38258 28512
rect 38562 28500 38568 28552
rect 38620 28540 38626 28552
rect 38841 28543 38899 28549
rect 38841 28540 38853 28543
rect 38620 28512 38853 28540
rect 38620 28500 38626 28512
rect 38841 28509 38853 28512
rect 38887 28509 38899 28543
rect 38841 28503 38899 28509
rect 39942 28500 39948 28552
rect 40000 28540 40006 28552
rect 40037 28543 40095 28549
rect 40037 28540 40049 28543
rect 40000 28512 40049 28540
rect 40000 28500 40006 28512
rect 40037 28509 40049 28512
rect 40083 28509 40095 28543
rect 40037 28503 40095 28509
rect 40126 28500 40132 28552
rect 40184 28540 40190 28552
rect 40184 28512 40229 28540
rect 40184 28500 40190 28512
rect 41138 28500 41144 28552
rect 41196 28540 41202 28552
rect 41524 28549 41552 28580
rect 42702 28568 42708 28580
rect 42760 28568 42766 28620
rect 41233 28543 41291 28549
rect 41233 28540 41245 28543
rect 41196 28512 41245 28540
rect 41196 28500 41202 28512
rect 41233 28509 41245 28512
rect 41279 28509 41291 28543
rect 41524 28543 41593 28549
rect 41524 28512 41547 28543
rect 41233 28503 41291 28509
rect 41535 28509 41547 28512
rect 41581 28509 41593 28543
rect 41535 28503 41593 28509
rect 41693 28543 41751 28549
rect 41693 28509 41705 28543
rect 41739 28509 41751 28543
rect 41693 28503 41751 28509
rect 31662 28432 31668 28484
rect 31720 28432 31726 28484
rect 32309 28475 32367 28481
rect 32309 28441 32321 28475
rect 32355 28472 32367 28475
rect 33778 28472 33784 28484
rect 32355 28444 33784 28472
rect 32355 28441 32367 28444
rect 32309 28435 32367 28441
rect 33778 28432 33784 28444
rect 33836 28432 33842 28484
rect 33134 28404 33140 28416
rect 33095 28376 33140 28404
rect 33134 28364 33140 28376
rect 33192 28364 33198 28416
rect 33689 28407 33747 28413
rect 33689 28373 33701 28407
rect 33735 28404 33747 28407
rect 35710 28404 35716 28416
rect 33735 28376 35716 28404
rect 33735 28373 33747 28376
rect 33689 28367 33747 28373
rect 35710 28364 35716 28376
rect 35768 28364 35774 28416
rect 35912 28404 35940 28500
rect 36078 28472 36084 28484
rect 36039 28444 36084 28472
rect 36078 28432 36084 28444
rect 36136 28432 36142 28484
rect 36219 28475 36277 28481
rect 36219 28441 36231 28475
rect 36265 28472 36277 28475
rect 37918 28472 37924 28484
rect 36265 28444 37924 28472
rect 36265 28441 36277 28444
rect 36219 28435 36277 28441
rect 37918 28432 37924 28444
rect 37976 28472 37982 28484
rect 37976 28444 38884 28472
rect 37976 28432 37982 28444
rect 37366 28404 37372 28416
rect 35912 28376 37372 28404
rect 37366 28364 37372 28376
rect 37424 28364 37430 28416
rect 38381 28407 38439 28413
rect 38381 28373 38393 28407
rect 38427 28404 38439 28407
rect 38654 28404 38660 28416
rect 38427 28376 38660 28404
rect 38427 28373 38439 28376
rect 38381 28367 38439 28373
rect 38654 28364 38660 28376
rect 38712 28364 38718 28416
rect 38856 28413 38884 28444
rect 38930 28432 38936 28484
rect 38988 28472 38994 28484
rect 39117 28475 39175 28481
rect 38988 28444 39033 28472
rect 38988 28432 38994 28444
rect 39117 28441 39129 28475
rect 39163 28472 39175 28475
rect 39206 28472 39212 28484
rect 39163 28444 39212 28472
rect 39163 28441 39175 28444
rect 39117 28435 39175 28441
rect 39206 28432 39212 28444
rect 39264 28432 39270 28484
rect 40862 28432 40868 28484
rect 40920 28472 40926 28484
rect 41325 28475 41383 28481
rect 41325 28472 41337 28475
rect 40920 28444 41337 28472
rect 40920 28432 40926 28444
rect 41325 28441 41337 28444
rect 41371 28441 41383 28475
rect 41325 28435 41383 28441
rect 41414 28432 41420 28484
rect 41472 28472 41478 28484
rect 41708 28472 41736 28503
rect 41782 28500 41788 28552
rect 41840 28540 41846 28552
rect 42337 28543 42395 28549
rect 42337 28540 42349 28543
rect 41840 28512 42349 28540
rect 41840 28500 41846 28512
rect 42337 28509 42349 28512
rect 42383 28509 42395 28543
rect 42337 28503 42395 28509
rect 41874 28472 41880 28484
rect 41472 28444 41517 28472
rect 41708 28444 41880 28472
rect 41472 28432 41478 28444
rect 41874 28432 41880 28444
rect 41932 28432 41938 28484
rect 42812 28472 42840 28648
rect 43254 28540 43260 28552
rect 43215 28512 43260 28540
rect 43254 28500 43260 28512
rect 43312 28500 43318 28552
rect 43364 28540 43392 28716
rect 45186 28704 45192 28716
rect 45244 28704 45250 28756
rect 45278 28704 45284 28756
rect 45336 28744 45342 28756
rect 47670 28744 47676 28756
rect 45336 28716 47676 28744
rect 45336 28704 45342 28716
rect 47670 28704 47676 28716
rect 47728 28744 47734 28756
rect 48225 28747 48283 28753
rect 48225 28744 48237 28747
rect 47728 28716 48237 28744
rect 47728 28704 47734 28716
rect 48225 28713 48237 28716
rect 48271 28713 48283 28747
rect 49326 28744 49332 28756
rect 48225 28707 48283 28713
rect 48332 28716 49332 28744
rect 44726 28676 44732 28688
rect 44008 28648 44732 28676
rect 44008 28617 44036 28648
rect 44726 28636 44732 28648
rect 44784 28676 44790 28688
rect 47302 28676 47308 28688
rect 44784 28648 47308 28676
rect 44784 28636 44790 28648
rect 47302 28636 47308 28648
rect 47360 28676 47366 28688
rect 48130 28676 48136 28688
rect 47360 28648 48136 28676
rect 47360 28636 47366 28648
rect 48130 28636 48136 28648
rect 48188 28676 48194 28688
rect 48332 28676 48360 28716
rect 49326 28704 49332 28716
rect 49384 28704 49390 28756
rect 49694 28704 49700 28756
rect 49752 28744 49758 28756
rect 50341 28747 50399 28753
rect 50341 28744 50353 28747
rect 49752 28716 50353 28744
rect 49752 28704 49758 28716
rect 50341 28713 50353 28716
rect 50387 28713 50399 28747
rect 50341 28707 50399 28713
rect 50540 28716 50752 28744
rect 48188 28648 48360 28676
rect 48188 28636 48194 28648
rect 48866 28636 48872 28688
rect 48924 28676 48930 28688
rect 50430 28676 50436 28688
rect 48924 28648 50436 28676
rect 48924 28636 48930 28648
rect 50430 28636 50436 28648
rect 50488 28636 50494 28688
rect 43993 28611 44051 28617
rect 43993 28577 44005 28611
rect 44039 28577 44051 28611
rect 43993 28571 44051 28577
rect 45186 28568 45192 28620
rect 45244 28608 45250 28620
rect 46842 28608 46848 28620
rect 45244 28580 45600 28608
rect 45244 28568 45250 28580
rect 45572 28549 45600 28580
rect 46400 28580 46848 28608
rect 44177 28543 44235 28549
rect 44177 28540 44189 28543
rect 43364 28512 44189 28540
rect 44177 28509 44189 28512
rect 44223 28540 44235 28543
rect 45327 28543 45385 28549
rect 45327 28540 45339 28543
rect 44223 28512 45339 28540
rect 44223 28509 44235 28512
rect 44177 28503 44235 28509
rect 45327 28509 45339 28512
rect 45373 28509 45385 28543
rect 45327 28503 45385 28509
rect 45557 28543 45615 28549
rect 45557 28509 45569 28543
rect 45603 28509 45615 28543
rect 45557 28503 45615 28509
rect 45646 28500 45652 28552
rect 45704 28549 45710 28552
rect 45704 28543 45743 28549
rect 45731 28509 45743 28543
rect 45704 28503 45743 28509
rect 45704 28500 45710 28503
rect 45830 28500 45836 28552
rect 45888 28540 45894 28552
rect 46290 28540 46296 28552
rect 45888 28512 45933 28540
rect 46251 28512 46296 28540
rect 45888 28500 45894 28512
rect 46290 28500 46296 28512
rect 46348 28500 46354 28552
rect 46400 28549 46428 28580
rect 46842 28568 46848 28580
rect 46900 28568 46906 28620
rect 48590 28608 48596 28620
rect 47320 28580 48596 28608
rect 46385 28543 46443 28549
rect 46385 28509 46397 28543
rect 46431 28509 46443 28543
rect 46385 28503 46443 28509
rect 46569 28543 46627 28549
rect 46569 28509 46581 28543
rect 46615 28540 46627 28543
rect 46658 28540 46664 28552
rect 46615 28512 46664 28540
rect 46615 28509 46627 28512
rect 46569 28503 46627 28509
rect 46658 28500 46664 28512
rect 46716 28540 46722 28552
rect 47320 28540 47348 28580
rect 48590 28568 48596 28580
rect 48648 28568 48654 28620
rect 49142 28608 49148 28620
rect 49103 28580 49148 28608
rect 49142 28568 49148 28580
rect 49200 28568 49206 28620
rect 49329 28611 49387 28617
rect 49329 28577 49341 28611
rect 49375 28608 49387 28611
rect 50540 28608 50568 28716
rect 49375 28580 50568 28608
rect 50724 28608 50752 28716
rect 52454 28704 52460 28756
rect 52512 28744 52518 28756
rect 55585 28747 55643 28753
rect 55585 28744 55597 28747
rect 52512 28716 55597 28744
rect 52512 28704 52518 28716
rect 55585 28713 55597 28716
rect 55631 28744 55643 28747
rect 56045 28747 56103 28753
rect 56045 28744 56057 28747
rect 55631 28716 56057 28744
rect 55631 28713 55643 28716
rect 55585 28707 55643 28713
rect 56045 28713 56057 28716
rect 56091 28713 56103 28747
rect 56045 28707 56103 28713
rect 50798 28636 50804 28688
rect 50856 28676 50862 28688
rect 51629 28679 51687 28685
rect 51629 28676 51641 28679
rect 50856 28648 51641 28676
rect 50856 28636 50862 28648
rect 51629 28645 51641 28648
rect 51675 28645 51687 28679
rect 54386 28676 54392 28688
rect 54347 28648 54392 28676
rect 51629 28639 51687 28645
rect 54386 28636 54392 28648
rect 54444 28636 54450 28688
rect 57330 28636 57336 28688
rect 57388 28676 57394 28688
rect 57388 28648 57928 28676
rect 57388 28636 57394 28648
rect 54846 28608 54852 28620
rect 50724 28580 51212 28608
rect 54807 28580 54852 28608
rect 49375 28577 49387 28580
rect 49329 28571 49387 28577
rect 47486 28540 47492 28552
rect 46716 28512 47348 28540
rect 47399 28512 47492 28540
rect 46716 28500 46722 28512
rect 47486 28500 47492 28512
rect 47544 28500 47550 28552
rect 47581 28543 47639 28549
rect 47581 28509 47593 28543
rect 47627 28540 47639 28543
rect 47670 28540 47676 28552
rect 47627 28512 47676 28540
rect 47627 28509 47639 28512
rect 47581 28503 47639 28509
rect 47670 28500 47676 28512
rect 47728 28500 47734 28552
rect 48222 28500 48228 28552
rect 48280 28540 48286 28552
rect 48409 28543 48467 28549
rect 48280 28512 48325 28540
rect 48280 28500 48286 28512
rect 48409 28509 48421 28543
rect 48455 28509 48467 28543
rect 49050 28540 49056 28552
rect 49011 28512 49056 28540
rect 48409 28503 48467 28509
rect 44085 28475 44143 28481
rect 44085 28472 44097 28475
rect 42812 28444 44097 28472
rect 44085 28441 44097 28444
rect 44131 28472 44143 28475
rect 45186 28472 45192 28484
rect 44131 28444 45192 28472
rect 44131 28441 44143 28444
rect 44085 28435 44143 28441
rect 45186 28432 45192 28444
rect 45244 28432 45250 28484
rect 45465 28475 45523 28481
rect 45465 28441 45477 28475
rect 45511 28472 45523 28475
rect 47302 28472 47308 28484
rect 45511 28444 47308 28472
rect 45511 28441 45523 28444
rect 45465 28435 45523 28441
rect 47302 28432 47308 28444
rect 47360 28432 47366 28484
rect 47504 28472 47532 28500
rect 48424 28472 48452 28503
rect 49050 28500 49056 28512
rect 49108 28500 49114 28552
rect 49418 28540 49424 28552
rect 49379 28512 49424 28540
rect 49418 28500 49424 28512
rect 49476 28500 49482 28552
rect 50338 28540 50344 28552
rect 50299 28512 50344 28540
rect 50338 28500 50344 28512
rect 50396 28500 50402 28552
rect 50522 28540 50528 28552
rect 50483 28512 50528 28540
rect 50522 28500 50528 28512
rect 50580 28500 50586 28552
rect 50614 28500 50620 28552
rect 50672 28540 50678 28552
rect 51184 28549 51212 28580
rect 54846 28568 54852 28580
rect 54904 28568 54910 28620
rect 57514 28568 57520 28620
rect 57572 28608 57578 28620
rect 57900 28617 57928 28648
rect 57793 28611 57851 28617
rect 57793 28608 57805 28611
rect 57572 28580 57805 28608
rect 57572 28568 57578 28580
rect 57793 28577 57805 28580
rect 57839 28577 57851 28611
rect 57793 28571 57851 28577
rect 57885 28611 57943 28617
rect 57885 28577 57897 28611
rect 57931 28577 57943 28611
rect 57885 28571 57943 28577
rect 50985 28543 51043 28549
rect 50985 28540 50997 28543
rect 50672 28512 50997 28540
rect 50672 28500 50678 28512
rect 50985 28509 50997 28512
rect 51031 28509 51043 28543
rect 50985 28503 51043 28509
rect 51169 28543 51227 28549
rect 51169 28509 51181 28543
rect 51215 28540 51227 28543
rect 51534 28540 51540 28552
rect 51215 28512 51540 28540
rect 51215 28509 51227 28512
rect 51169 28503 51227 28509
rect 51534 28500 51540 28512
rect 51592 28500 51598 28552
rect 52270 28540 52276 28552
rect 52231 28512 52276 28540
rect 52270 28500 52276 28512
rect 52328 28500 52334 28552
rect 53374 28540 53380 28552
rect 53335 28512 53380 28540
rect 53374 28500 53380 28512
rect 53432 28500 53438 28552
rect 53466 28500 53472 28552
rect 53524 28540 53530 28552
rect 53524 28512 53569 28540
rect 53524 28500 53530 28512
rect 53650 28500 53656 28552
rect 53708 28549 53714 28552
rect 53708 28543 53737 28549
rect 53725 28509 53737 28543
rect 53708 28503 53737 28509
rect 53837 28543 53895 28549
rect 53837 28509 53849 28543
rect 53883 28540 53895 28543
rect 54110 28540 54116 28552
rect 53883 28512 54116 28540
rect 53883 28509 53895 28512
rect 53837 28503 53895 28509
rect 53708 28500 53714 28503
rect 54110 28500 54116 28512
rect 54168 28500 54174 28552
rect 54754 28540 54760 28552
rect 54715 28512 54760 28540
rect 54754 28500 54760 28512
rect 54812 28500 54818 28552
rect 57238 28500 57244 28552
rect 57296 28540 57302 28552
rect 57701 28543 57759 28549
rect 57701 28540 57713 28543
rect 57296 28512 57713 28540
rect 57296 28500 57302 28512
rect 57701 28509 57713 28512
rect 57747 28509 57759 28543
rect 57701 28503 57759 28509
rect 52365 28475 52423 28481
rect 52365 28472 52377 28475
rect 47504 28444 52377 28472
rect 52365 28441 52377 28444
rect 52411 28472 52423 28475
rect 53561 28475 53619 28481
rect 53561 28472 53573 28475
rect 52411 28444 53573 28472
rect 52411 28441 52423 28444
rect 52365 28435 52423 28441
rect 53561 28441 53573 28444
rect 53607 28472 53619 28475
rect 54018 28472 54024 28484
rect 53607 28444 54024 28472
rect 53607 28441 53619 28444
rect 53561 28435 53619 28441
rect 54018 28432 54024 28444
rect 54076 28432 54082 28484
rect 38841 28407 38899 28413
rect 38841 28373 38853 28407
rect 38887 28373 38899 28407
rect 41046 28404 41052 28416
rect 41007 28376 41052 28404
rect 38841 28367 38899 28373
rect 41046 28364 41052 28376
rect 41104 28364 41110 28416
rect 42150 28404 42156 28416
rect 42111 28376 42156 28404
rect 42150 28364 42156 28376
rect 42208 28364 42214 28416
rect 42242 28364 42248 28416
rect 42300 28404 42306 28416
rect 43165 28407 43223 28413
rect 43165 28404 43177 28407
rect 42300 28376 43177 28404
rect 42300 28364 42306 28376
rect 43165 28373 43177 28376
rect 43211 28404 43223 28407
rect 44266 28404 44272 28416
rect 43211 28376 44272 28404
rect 43211 28373 43223 28376
rect 43165 28367 43223 28373
rect 44266 28364 44272 28376
rect 44324 28364 44330 28416
rect 44545 28407 44603 28413
rect 44545 28373 44557 28407
rect 44591 28404 44603 28407
rect 46106 28404 46112 28416
rect 44591 28376 46112 28404
rect 44591 28373 44603 28376
rect 44545 28367 44603 28373
rect 46106 28364 46112 28376
rect 46164 28364 46170 28416
rect 46750 28404 46756 28416
rect 46711 28376 46756 28404
rect 46750 28364 46756 28376
rect 46808 28364 46814 28416
rect 47320 28404 47348 28432
rect 47765 28407 47823 28413
rect 47765 28404 47777 28407
rect 47320 28376 47777 28404
rect 47765 28373 47777 28376
rect 47811 28404 47823 28407
rect 47854 28404 47860 28416
rect 47811 28376 47860 28404
rect 47811 28373 47823 28376
rect 47765 28367 47823 28373
rect 47854 28364 47860 28376
rect 47912 28364 47918 28416
rect 49053 28407 49111 28413
rect 49053 28373 49065 28407
rect 49099 28404 49111 28407
rect 49326 28404 49332 28416
rect 49099 28376 49332 28404
rect 49099 28373 49111 28376
rect 49053 28367 49111 28373
rect 49326 28364 49332 28376
rect 49384 28364 49390 28416
rect 51074 28404 51080 28416
rect 51035 28376 51080 28404
rect 51074 28364 51080 28376
rect 51132 28364 51138 28416
rect 53193 28407 53251 28413
rect 53193 28373 53205 28407
rect 53239 28404 53251 28407
rect 53926 28404 53932 28416
rect 53239 28376 53932 28404
rect 53239 28373 53251 28376
rect 53193 28367 53251 28373
rect 53926 28364 53932 28376
rect 53984 28364 53990 28416
rect 56594 28404 56600 28416
rect 56555 28376 56600 28404
rect 56594 28364 56600 28376
rect 56652 28364 56658 28416
rect 57238 28364 57244 28416
rect 57296 28404 57302 28416
rect 57333 28407 57391 28413
rect 57333 28404 57345 28407
rect 57296 28376 57345 28404
rect 57296 28364 57302 28376
rect 57333 28373 57345 28376
rect 57379 28373 57391 28407
rect 57333 28367 57391 28373
rect 1104 28314 58880 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 58880 28314
rect 1104 28240 58880 28262
rect 37366 28160 37372 28212
rect 37424 28200 37430 28212
rect 37553 28203 37611 28209
rect 37553 28200 37565 28203
rect 37424 28172 37565 28200
rect 37424 28160 37430 28172
rect 37553 28169 37565 28172
rect 37599 28169 37611 28203
rect 38286 28200 38292 28212
rect 38247 28172 38292 28200
rect 37553 28163 37611 28169
rect 38286 28160 38292 28172
rect 38344 28160 38350 28212
rect 40129 28203 40187 28209
rect 40129 28169 40141 28203
rect 40175 28200 40187 28203
rect 40310 28200 40316 28212
rect 40175 28172 40316 28200
rect 40175 28169 40187 28172
rect 40129 28163 40187 28169
rect 40310 28160 40316 28172
rect 40368 28160 40374 28212
rect 41417 28203 41475 28209
rect 41417 28169 41429 28203
rect 41463 28200 41475 28203
rect 41782 28200 41788 28212
rect 41463 28172 41552 28200
rect 41743 28172 41788 28200
rect 41463 28169 41475 28172
rect 41417 28163 41475 28169
rect 33134 28092 33140 28144
rect 33192 28092 33198 28144
rect 34330 28132 34336 28144
rect 34291 28104 34336 28132
rect 34330 28092 34336 28104
rect 34388 28092 34394 28144
rect 34514 28092 34520 28144
rect 34572 28132 34578 28144
rect 34793 28135 34851 28141
rect 34793 28132 34805 28135
rect 34572 28104 34805 28132
rect 34572 28092 34578 28104
rect 34793 28101 34805 28104
rect 34839 28101 34851 28135
rect 34793 28095 34851 28101
rect 37550 28024 37556 28076
rect 37608 28064 37614 28076
rect 37737 28067 37795 28073
rect 37737 28064 37749 28067
rect 37608 28036 37749 28064
rect 37608 28024 37614 28036
rect 37737 28033 37749 28036
rect 37783 28064 37795 28067
rect 38841 28067 38899 28073
rect 38841 28064 38853 28067
rect 37783 28036 38853 28064
rect 37783 28033 37795 28036
rect 37737 28027 37795 28033
rect 38841 28033 38853 28036
rect 38887 28064 38899 28067
rect 39206 28064 39212 28076
rect 38887 28036 39212 28064
rect 38887 28033 38899 28036
rect 38841 28027 38899 28033
rect 39206 28024 39212 28036
rect 39264 28024 39270 28076
rect 39761 28067 39819 28073
rect 39761 28033 39773 28067
rect 39807 28033 39819 28067
rect 41524 28064 41552 28172
rect 41782 28160 41788 28172
rect 41840 28160 41846 28212
rect 41874 28160 41880 28212
rect 41932 28200 41938 28212
rect 43162 28200 43168 28212
rect 41932 28172 43168 28200
rect 41932 28160 41938 28172
rect 43162 28160 43168 28172
rect 43220 28200 43226 28212
rect 43714 28200 43720 28212
rect 43220 28172 43720 28200
rect 43220 28160 43226 28172
rect 43714 28160 43720 28172
rect 43772 28160 43778 28212
rect 44174 28160 44180 28212
rect 44232 28200 44238 28212
rect 45373 28203 45431 28209
rect 45373 28200 45385 28203
rect 44232 28172 45385 28200
rect 44232 28160 44238 28172
rect 45373 28169 45385 28172
rect 45419 28200 45431 28203
rect 45462 28200 45468 28212
rect 45419 28172 45468 28200
rect 45419 28169 45431 28172
rect 45373 28163 45431 28169
rect 45462 28160 45468 28172
rect 45520 28160 45526 28212
rect 45741 28203 45799 28209
rect 45741 28169 45753 28203
rect 45787 28200 45799 28203
rect 46290 28200 46296 28212
rect 45787 28172 46296 28200
rect 45787 28169 45799 28172
rect 45741 28163 45799 28169
rect 46290 28160 46296 28172
rect 46348 28160 46354 28212
rect 47118 28160 47124 28212
rect 47176 28200 47182 28212
rect 49602 28200 49608 28212
rect 47176 28172 49608 28200
rect 47176 28160 47182 28172
rect 49602 28160 49608 28172
rect 49660 28160 49666 28212
rect 49694 28160 49700 28212
rect 49752 28200 49758 28212
rect 50522 28200 50528 28212
rect 49752 28172 50528 28200
rect 49752 28160 49758 28172
rect 50522 28160 50528 28172
rect 50580 28200 50586 28212
rect 51994 28200 52000 28212
rect 50580 28172 51074 28200
rect 51955 28172 52000 28200
rect 50580 28160 50586 28172
rect 45278 28132 45284 28144
rect 44192 28104 45284 28132
rect 42242 28064 42248 28076
rect 41524 28036 42248 28064
rect 39761 28027 39819 28033
rect 32306 27996 32312 28008
rect 32267 27968 32312 27996
rect 32306 27956 32312 27968
rect 32364 27956 32370 28008
rect 32582 27996 32588 28008
rect 32543 27968 32588 27996
rect 32582 27956 32588 27968
rect 32640 27956 32646 28008
rect 38378 27956 38384 28008
rect 38436 27996 38442 28008
rect 38562 27996 38568 28008
rect 38436 27968 38568 27996
rect 38436 27956 38442 27968
rect 38562 27956 38568 27968
rect 38620 27996 38626 28008
rect 39482 27996 39488 28008
rect 38620 27968 39488 27996
rect 38620 27956 38626 27968
rect 39482 27956 39488 27968
rect 39540 27956 39546 28008
rect 37274 27888 37280 27940
rect 37332 27928 37338 27940
rect 39776 27928 39804 28027
rect 42242 28024 42248 28036
rect 42300 28024 42306 28076
rect 42518 28024 42524 28076
rect 42576 28064 42582 28076
rect 42613 28067 42671 28073
rect 42613 28064 42625 28067
rect 42576 28036 42625 28064
rect 42576 28024 42582 28036
rect 42613 28033 42625 28036
rect 42659 28033 42671 28067
rect 42613 28027 42671 28033
rect 43901 28067 43959 28073
rect 43901 28033 43913 28067
rect 43947 28033 43959 28067
rect 43901 28027 43959 28033
rect 39853 27999 39911 28005
rect 39853 27965 39865 27999
rect 39899 27996 39911 27999
rect 40126 27996 40132 28008
rect 39899 27968 40132 27996
rect 39899 27965 39911 27968
rect 39853 27959 39911 27965
rect 37332 27900 39804 27928
rect 37332 27888 37338 27900
rect 31754 27820 31760 27872
rect 31812 27860 31818 27872
rect 31812 27832 31857 27860
rect 31812 27820 31818 27832
rect 32950 27820 32956 27872
rect 33008 27860 33014 27872
rect 36081 27863 36139 27869
rect 36081 27860 36093 27863
rect 33008 27832 36093 27860
rect 33008 27820 33014 27832
rect 36081 27829 36093 27832
rect 36127 27829 36139 27863
rect 36081 27823 36139 27829
rect 38749 27863 38807 27869
rect 38749 27829 38761 27863
rect 38795 27860 38807 27863
rect 39022 27860 39028 27872
rect 38795 27832 39028 27860
rect 38795 27829 38807 27832
rect 38749 27823 38807 27829
rect 39022 27820 39028 27832
rect 39080 27820 39086 27872
rect 39482 27820 39488 27872
rect 39540 27860 39546 27872
rect 39868 27860 39896 27959
rect 40126 27956 40132 27968
rect 40184 27956 40190 28008
rect 41233 27999 41291 28005
rect 41233 27965 41245 27999
rect 41279 27965 41291 27999
rect 41233 27959 41291 27965
rect 41325 27999 41383 28005
rect 41325 27965 41337 27999
rect 41371 27996 41383 27999
rect 41966 27996 41972 28008
rect 41371 27968 41972 27996
rect 41371 27965 41383 27968
rect 41325 27959 41383 27965
rect 41248 27928 41276 27959
rect 41966 27956 41972 27968
rect 42024 27996 42030 28008
rect 43257 27999 43315 28005
rect 43257 27996 43269 27999
rect 42024 27968 43269 27996
rect 42024 27956 42030 27968
rect 43257 27965 43269 27968
rect 43303 27996 43315 27999
rect 43806 27996 43812 28008
rect 43303 27968 43812 27996
rect 43303 27965 43315 27968
rect 43257 27959 43315 27965
rect 43806 27956 43812 27968
rect 43864 27956 43870 28008
rect 43916 27996 43944 28027
rect 43990 28024 43996 28076
rect 44048 28064 44054 28076
rect 44192 28073 44220 28104
rect 45278 28092 45284 28104
rect 45336 28092 45342 28144
rect 46845 28135 46903 28141
rect 46845 28101 46857 28135
rect 46891 28132 46903 28135
rect 46891 28104 49464 28132
rect 46891 28101 46903 28104
rect 46845 28095 46903 28101
rect 44177 28067 44235 28073
rect 44048 28036 44093 28064
rect 44048 28024 44054 28036
rect 44177 28033 44189 28067
rect 44223 28033 44235 28067
rect 44177 28027 44235 28033
rect 44266 28024 44272 28076
rect 44324 28064 44330 28076
rect 44407 28067 44465 28073
rect 44324 28036 44369 28064
rect 44324 28024 44330 28036
rect 44407 28033 44419 28067
rect 44453 28064 44465 28067
rect 45646 28064 45652 28076
rect 44453 28036 45652 28064
rect 44453 28033 44465 28036
rect 44407 28027 44465 28033
rect 45646 28024 45652 28036
rect 45704 28024 45710 28076
rect 46201 28067 46259 28073
rect 46201 28033 46213 28067
rect 46247 28033 46259 28067
rect 46382 28064 46388 28076
rect 46343 28036 46388 28064
rect 46201 28027 46259 28033
rect 45002 27996 45008 28008
rect 43916 27968 45008 27996
rect 45002 27956 45008 27968
rect 45060 27956 45066 28008
rect 45189 27999 45247 28005
rect 45189 27965 45201 27999
rect 45235 27965 45247 27999
rect 45189 27959 45247 27965
rect 41414 27928 41420 27940
rect 41248 27900 41420 27928
rect 41414 27888 41420 27900
rect 41472 27888 41478 27940
rect 45204 27928 45232 27959
rect 45278 27956 45284 28008
rect 45336 27996 45342 28008
rect 45922 27996 45928 28008
rect 45336 27968 45928 27996
rect 45336 27956 45342 27968
rect 45922 27956 45928 27968
rect 45980 27956 45986 28008
rect 46216 27996 46244 28027
rect 46382 28024 46388 28036
rect 46440 28024 46446 28076
rect 46474 28024 46480 28076
rect 46532 28064 46538 28076
rect 46658 28073 46664 28076
rect 46615 28067 46664 28073
rect 46532 28036 46577 28064
rect 46532 28024 46538 28036
rect 46615 28033 46627 28067
rect 46661 28033 46664 28067
rect 46615 28027 46664 28033
rect 46658 28024 46664 28027
rect 46716 28024 46722 28076
rect 47765 28067 47823 28073
rect 47765 28033 47777 28067
rect 47811 28064 47823 28067
rect 47854 28064 47860 28076
rect 47811 28036 47860 28064
rect 47811 28033 47823 28036
rect 47765 28027 47823 28033
rect 47854 28024 47860 28036
rect 47912 28024 47918 28076
rect 47949 28067 48007 28073
rect 47949 28033 47961 28067
rect 47995 28064 48007 28067
rect 48038 28064 48044 28076
rect 47995 28036 48044 28064
rect 47995 28033 48007 28036
rect 47949 28027 48007 28033
rect 48038 28024 48044 28036
rect 48096 28024 48102 28076
rect 48774 28064 48780 28076
rect 48735 28036 48780 28064
rect 48774 28024 48780 28036
rect 48832 28024 48838 28076
rect 48958 28064 48964 28076
rect 48919 28036 48964 28064
rect 48958 28024 48964 28036
rect 49016 28024 49022 28076
rect 49436 28064 49464 28104
rect 50338 28092 50344 28144
rect 50396 28132 50402 28144
rect 51046 28132 51074 28172
rect 51994 28160 52000 28172
rect 52052 28160 52058 28212
rect 53374 28160 53380 28212
rect 53432 28200 53438 28212
rect 53653 28203 53711 28209
rect 53653 28200 53665 28203
rect 53432 28172 53665 28200
rect 53432 28160 53438 28172
rect 53653 28169 53665 28172
rect 53699 28169 53711 28203
rect 53653 28163 53711 28169
rect 54297 28203 54355 28209
rect 54297 28169 54309 28203
rect 54343 28200 54355 28203
rect 55214 28200 55220 28212
rect 54343 28172 55220 28200
rect 54343 28169 54355 28172
rect 54297 28163 54355 28169
rect 55214 28160 55220 28172
rect 55272 28160 55278 28212
rect 52270 28132 52276 28144
rect 50396 28104 50844 28132
rect 51046 28104 52276 28132
rect 50396 28092 50402 28104
rect 49973 28067 50031 28073
rect 49973 28064 49985 28067
rect 49436 28036 49985 28064
rect 49973 28033 49985 28036
rect 50019 28033 50031 28067
rect 49973 28027 50031 28033
rect 50065 28067 50123 28073
rect 50065 28033 50077 28067
rect 50111 28064 50123 28067
rect 50614 28064 50620 28076
rect 50111 28036 50620 28064
rect 50111 28033 50123 28036
rect 50065 28027 50123 28033
rect 50614 28024 50620 28036
rect 50672 28024 50678 28076
rect 50816 28064 50844 28104
rect 52270 28092 52276 28104
rect 52328 28092 52334 28144
rect 52822 28092 52828 28144
rect 52880 28132 52886 28144
rect 53285 28135 53343 28141
rect 53285 28132 53297 28135
rect 52880 28104 53297 28132
rect 52880 28092 52886 28104
rect 53285 28101 53297 28104
rect 53331 28101 53343 28135
rect 53285 28095 53343 28101
rect 53469 28135 53527 28141
rect 53469 28101 53481 28135
rect 53515 28132 53527 28135
rect 53558 28132 53564 28144
rect 53515 28104 53564 28132
rect 53515 28101 53527 28104
rect 53469 28095 53527 28101
rect 53558 28092 53564 28104
rect 53616 28092 53622 28144
rect 54018 28092 54024 28144
rect 54076 28132 54082 28144
rect 54113 28135 54171 28141
rect 54113 28132 54125 28135
rect 54076 28104 54125 28132
rect 54076 28092 54082 28104
rect 54113 28101 54125 28104
rect 54159 28101 54171 28135
rect 54113 28095 54171 28101
rect 51077 28067 51135 28073
rect 51077 28064 51089 28067
rect 50816 28036 51089 28064
rect 51077 28033 51089 28036
rect 51123 28033 51135 28067
rect 51350 28064 51356 28076
rect 51311 28036 51356 28064
rect 51077 28027 51135 28033
rect 51350 28024 51356 28036
rect 51408 28024 51414 28076
rect 51534 28064 51540 28076
rect 51495 28036 51540 28064
rect 51534 28024 51540 28036
rect 51592 28024 51598 28076
rect 54386 28024 54392 28076
rect 54444 28064 54450 28076
rect 55232 28064 55260 28160
rect 55493 28067 55551 28073
rect 55493 28064 55505 28067
rect 54444 28036 54489 28064
rect 55232 28036 55505 28064
rect 54444 28024 54450 28036
rect 55493 28033 55505 28036
rect 55539 28033 55551 28067
rect 57146 28064 57152 28076
rect 57107 28036 57152 28064
rect 55493 28027 55551 28033
rect 57146 28024 57152 28036
rect 57204 28024 57210 28076
rect 58342 28064 58348 28076
rect 58303 28036 58348 28064
rect 58342 28024 58348 28036
rect 58400 28024 58406 28076
rect 49602 27996 49608 28008
rect 46216 27968 49608 27996
rect 49602 27956 49608 27968
rect 49660 27956 49666 28008
rect 50157 27999 50215 28005
rect 50157 27996 50169 27999
rect 49712 27968 50169 27996
rect 49145 27931 49203 27937
rect 45204 27900 45508 27928
rect 39540 27832 39896 27860
rect 39945 27863 40003 27869
rect 39540 27820 39546 27832
rect 39945 27829 39957 27863
rect 39991 27860 40003 27863
rect 40126 27860 40132 27872
rect 39991 27832 40132 27860
rect 39991 27829 40003 27832
rect 39945 27823 40003 27829
rect 40126 27820 40132 27832
rect 40184 27820 40190 27872
rect 42705 27863 42763 27869
rect 42705 27829 42717 27863
rect 42751 27860 42763 27863
rect 42978 27860 42984 27872
rect 42751 27832 42984 27860
rect 42751 27829 42763 27832
rect 42705 27823 42763 27829
rect 42978 27820 42984 27832
rect 43036 27820 43042 27872
rect 44545 27863 44603 27869
rect 44545 27829 44557 27863
rect 44591 27860 44603 27863
rect 45370 27860 45376 27872
rect 44591 27832 45376 27860
rect 44591 27829 44603 27832
rect 44545 27823 44603 27829
rect 45370 27820 45376 27832
rect 45428 27820 45434 27872
rect 45480 27860 45508 27900
rect 49145 27897 49157 27931
rect 49191 27928 49203 27931
rect 49712 27928 49740 27968
rect 50157 27965 50169 27968
rect 50203 27965 50215 27999
rect 50157 27959 50215 27965
rect 50246 27956 50252 28008
rect 50304 27996 50310 28008
rect 50304 27968 50349 27996
rect 50304 27956 50310 27968
rect 50430 27956 50436 28008
rect 50488 27996 50494 28008
rect 55582 27996 55588 28008
rect 50488 27968 55444 27996
rect 55543 27968 55588 27996
rect 50488 27956 50494 27968
rect 54110 27928 54116 27940
rect 49191 27900 49740 27928
rect 54071 27900 54116 27928
rect 49191 27897 49203 27900
rect 49145 27891 49203 27897
rect 54110 27888 54116 27900
rect 54168 27888 54174 27940
rect 55416 27928 55444 27968
rect 55582 27956 55588 27968
rect 55640 27956 55646 28008
rect 57238 27996 57244 28008
rect 57199 27968 57244 27996
rect 57238 27956 57244 27968
rect 57296 27956 57302 28008
rect 58066 27996 58072 28008
rect 58027 27968 58072 27996
rect 58066 27956 58072 27968
rect 58124 27956 58130 28008
rect 57330 27928 57336 27940
rect 55416 27900 57336 27928
rect 57330 27888 57336 27900
rect 57388 27888 57394 27940
rect 57517 27931 57575 27937
rect 57517 27897 57529 27931
rect 57563 27928 57575 27931
rect 58253 27931 58311 27937
rect 58253 27928 58265 27931
rect 57563 27900 58265 27928
rect 57563 27897 57575 27900
rect 57517 27891 57575 27897
rect 58253 27897 58265 27900
rect 58299 27897 58311 27931
rect 58253 27891 58311 27897
rect 47118 27860 47124 27872
rect 45480 27832 47124 27860
rect 47118 27820 47124 27832
rect 47176 27820 47182 27872
rect 47857 27863 47915 27869
rect 47857 27829 47869 27863
rect 47903 27860 47915 27863
rect 47946 27860 47952 27872
rect 47903 27832 47952 27860
rect 47903 27829 47915 27832
rect 47857 27823 47915 27829
rect 47946 27820 47952 27832
rect 48004 27820 48010 27872
rect 48961 27863 49019 27869
rect 48961 27829 48973 27863
rect 49007 27860 49019 27863
rect 49786 27860 49792 27872
rect 49007 27832 49792 27860
rect 49007 27829 49019 27832
rect 48961 27823 49019 27829
rect 49786 27820 49792 27832
rect 49844 27820 49850 27872
rect 50433 27863 50491 27869
rect 50433 27829 50445 27863
rect 50479 27860 50491 27863
rect 50522 27860 50528 27872
rect 50479 27832 50528 27860
rect 50479 27829 50491 27832
rect 50433 27823 50491 27829
rect 50522 27820 50528 27832
rect 50580 27820 50586 27872
rect 50893 27863 50951 27869
rect 50893 27829 50905 27863
rect 50939 27860 50951 27863
rect 51166 27860 51172 27872
rect 50939 27832 51172 27860
rect 50939 27829 50951 27832
rect 50893 27823 50951 27829
rect 51166 27820 51172 27832
rect 51224 27820 51230 27872
rect 55858 27860 55864 27872
rect 55819 27832 55864 27860
rect 55858 27820 55864 27832
rect 55916 27820 55922 27872
rect 56318 27860 56324 27872
rect 56279 27832 56324 27860
rect 56318 27820 56324 27832
rect 56376 27820 56382 27872
rect 57698 27820 57704 27872
rect 57756 27860 57762 27872
rect 58161 27863 58219 27869
rect 58161 27860 58173 27863
rect 57756 27832 58173 27860
rect 57756 27820 57762 27832
rect 58161 27829 58173 27832
rect 58207 27829 58219 27863
rect 58161 27823 58219 27829
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 32582 27656 32588 27668
rect 32543 27628 32588 27656
rect 32582 27616 32588 27628
rect 32640 27616 32646 27668
rect 37093 27659 37151 27665
rect 37093 27625 37105 27659
rect 37139 27656 37151 27659
rect 37182 27656 37188 27668
rect 37139 27628 37188 27656
rect 37139 27625 37151 27628
rect 37093 27619 37151 27625
rect 37182 27616 37188 27628
rect 37240 27616 37246 27668
rect 38194 27616 38200 27668
rect 38252 27656 38258 27668
rect 38562 27656 38568 27668
rect 38252 27628 38568 27656
rect 38252 27616 38258 27628
rect 38562 27616 38568 27628
rect 38620 27616 38626 27668
rect 39942 27616 39948 27668
rect 40000 27656 40006 27668
rect 40037 27659 40095 27665
rect 40037 27656 40049 27659
rect 40000 27628 40049 27656
rect 40000 27616 40006 27628
rect 40037 27625 40049 27628
rect 40083 27656 40095 27659
rect 40126 27656 40132 27668
rect 40083 27628 40132 27656
rect 40083 27625 40095 27628
rect 40037 27619 40095 27625
rect 40126 27616 40132 27628
rect 40184 27616 40190 27668
rect 40862 27616 40868 27668
rect 40920 27656 40926 27668
rect 40957 27659 41015 27665
rect 40957 27656 40969 27659
rect 40920 27628 40969 27656
rect 40920 27616 40926 27628
rect 40957 27625 40969 27628
rect 41003 27625 41015 27659
rect 40957 27619 41015 27625
rect 41956 27659 42014 27665
rect 41956 27625 41968 27659
rect 42002 27656 42014 27659
rect 42150 27656 42156 27668
rect 42002 27628 42156 27656
rect 42002 27625 42014 27628
rect 41956 27619 42014 27625
rect 42150 27616 42156 27628
rect 42208 27616 42214 27668
rect 43254 27616 43260 27668
rect 43312 27656 43318 27668
rect 43441 27659 43499 27665
rect 43441 27656 43453 27659
rect 43312 27628 43453 27656
rect 43312 27616 43318 27628
rect 43441 27625 43453 27628
rect 43487 27625 43499 27659
rect 43441 27619 43499 27625
rect 44358 27616 44364 27668
rect 44416 27656 44422 27668
rect 45278 27656 45284 27668
rect 44416 27628 45284 27656
rect 44416 27616 44422 27628
rect 45278 27616 45284 27628
rect 45336 27616 45342 27668
rect 46382 27616 46388 27668
rect 46440 27656 46446 27668
rect 46569 27659 46627 27665
rect 46569 27656 46581 27659
rect 46440 27628 46581 27656
rect 46440 27616 46446 27628
rect 46569 27625 46581 27628
rect 46615 27625 46627 27659
rect 46569 27619 46627 27625
rect 47118 27616 47124 27668
rect 47176 27656 47182 27668
rect 47670 27656 47676 27668
rect 47176 27628 47676 27656
rect 47176 27616 47182 27628
rect 47670 27616 47676 27628
rect 47728 27656 47734 27668
rect 49878 27656 49884 27668
rect 47728 27628 49884 27656
rect 47728 27616 47734 27628
rect 35253 27591 35311 27597
rect 35253 27557 35265 27591
rect 35299 27557 35311 27591
rect 36630 27588 36636 27600
rect 35253 27551 35311 27557
rect 35728 27560 36636 27588
rect 35268 27520 35296 27551
rect 35728 27529 35756 27560
rect 36630 27548 36636 27560
rect 36688 27548 36694 27600
rect 37274 27588 37280 27600
rect 37235 27560 37280 27588
rect 37274 27548 37280 27560
rect 37332 27548 37338 27600
rect 32784 27492 35296 27520
rect 35713 27523 35771 27529
rect 32784 27461 32812 27492
rect 35713 27489 35725 27523
rect 35759 27489 35771 27523
rect 35713 27483 35771 27489
rect 35897 27523 35955 27529
rect 35897 27489 35909 27523
rect 35943 27520 35955 27523
rect 36262 27520 36268 27532
rect 35943 27492 36268 27520
rect 35943 27489 35955 27492
rect 35897 27483 35955 27489
rect 32769 27455 32827 27461
rect 32769 27421 32781 27455
rect 32815 27421 32827 27455
rect 33778 27452 33784 27464
rect 33739 27424 33784 27452
rect 32769 27415 32827 27421
rect 33778 27412 33784 27424
rect 33836 27412 33842 27464
rect 34606 27412 34612 27464
rect 34664 27452 34670 27464
rect 35621 27455 35679 27461
rect 35621 27452 35633 27455
rect 34664 27424 35633 27452
rect 34664 27412 34670 27424
rect 35621 27421 35633 27424
rect 35667 27421 35679 27455
rect 35621 27415 35679 27421
rect 34333 27387 34391 27393
rect 34333 27353 34345 27387
rect 34379 27384 34391 27387
rect 35728 27384 35756 27483
rect 36262 27480 36268 27492
rect 36320 27480 36326 27532
rect 38212 27520 38240 27616
rect 38746 27588 38752 27600
rect 38707 27560 38752 27588
rect 38746 27548 38752 27560
rect 38804 27548 38810 27600
rect 39485 27591 39543 27597
rect 39485 27557 39497 27591
rect 39531 27588 39543 27591
rect 39574 27588 39580 27600
rect 39531 27560 39580 27588
rect 39531 27557 39543 27560
rect 39485 27551 39543 27557
rect 39574 27548 39580 27560
rect 39632 27548 39638 27600
rect 40405 27591 40463 27597
rect 40405 27557 40417 27591
rect 40451 27588 40463 27591
rect 40586 27588 40592 27600
rect 40451 27560 40592 27588
rect 40451 27557 40463 27560
rect 40405 27551 40463 27557
rect 40586 27548 40592 27560
rect 40644 27548 40650 27600
rect 46842 27548 46848 27600
rect 46900 27588 46906 27600
rect 47489 27591 47547 27597
rect 47489 27588 47501 27591
rect 46900 27560 47501 27588
rect 46900 27548 46906 27560
rect 47489 27557 47501 27560
rect 47535 27557 47547 27591
rect 47489 27551 47547 27557
rect 36740 27492 38240 27520
rect 36740 27461 36768 27492
rect 39022 27480 39028 27532
rect 39080 27520 39086 27532
rect 41598 27520 41604 27532
rect 39080 27492 40080 27520
rect 39080 27480 39086 27492
rect 36725 27455 36783 27461
rect 36725 27421 36737 27455
rect 36771 27421 36783 27455
rect 36725 27415 36783 27421
rect 37093 27455 37151 27461
rect 37093 27421 37105 27455
rect 37139 27452 37151 27455
rect 38194 27452 38200 27464
rect 37139 27424 38200 27452
rect 37139 27421 37151 27424
rect 37093 27415 37151 27421
rect 38194 27412 38200 27424
rect 38252 27412 38258 27464
rect 38654 27412 38660 27464
rect 38712 27452 38718 27464
rect 39393 27455 39451 27461
rect 39393 27452 39405 27455
rect 38712 27424 39405 27452
rect 38712 27412 38718 27424
rect 39393 27421 39405 27424
rect 39439 27421 39451 27455
rect 39393 27415 39451 27421
rect 39482 27412 39488 27464
rect 39540 27452 39546 27464
rect 40052 27461 40080 27492
rect 41386 27492 41604 27520
rect 40037 27455 40095 27461
rect 39540 27424 39585 27452
rect 39540 27412 39546 27424
rect 40037 27421 40049 27455
rect 40083 27421 40095 27455
rect 40037 27415 40095 27421
rect 40221 27455 40279 27461
rect 40221 27421 40233 27455
rect 40267 27452 40279 27455
rect 40678 27452 40684 27464
rect 40267 27424 40684 27452
rect 40267 27421 40279 27424
rect 40221 27415 40279 27421
rect 40678 27412 40684 27424
rect 40736 27412 40742 27464
rect 41141 27455 41199 27461
rect 41141 27421 41153 27455
rect 41187 27452 41199 27455
rect 41386 27452 41414 27492
rect 41598 27480 41604 27492
rect 41656 27480 41662 27532
rect 41693 27523 41751 27529
rect 41693 27489 41705 27523
rect 41739 27520 41751 27523
rect 42702 27520 42708 27532
rect 41739 27492 42708 27520
rect 41739 27489 41751 27492
rect 41693 27483 41751 27489
rect 42702 27480 42708 27492
rect 42760 27480 42766 27532
rect 48038 27520 48044 27532
rect 47688 27492 48044 27520
rect 44082 27452 44088 27464
rect 41187 27424 41414 27452
rect 44043 27424 44088 27452
rect 41187 27421 41199 27424
rect 41141 27415 41199 27421
rect 44082 27412 44088 27424
rect 44140 27412 44146 27464
rect 45370 27452 45376 27464
rect 45331 27424 45376 27452
rect 45370 27412 45376 27424
rect 45428 27412 45434 27464
rect 45462 27412 45468 27464
rect 45520 27452 45526 27464
rect 45649 27455 45707 27461
rect 45649 27452 45661 27455
rect 45520 27424 45661 27452
rect 45520 27412 45526 27424
rect 45649 27421 45661 27424
rect 45695 27421 45707 27455
rect 46106 27452 46112 27464
rect 46067 27424 46112 27452
rect 45649 27415 45707 27421
rect 46106 27412 46112 27424
rect 46164 27412 46170 27464
rect 46385 27455 46443 27461
rect 46385 27421 46397 27455
rect 46431 27452 46443 27455
rect 46750 27452 46756 27464
rect 46431 27424 46756 27452
rect 46431 27421 46443 27424
rect 46385 27415 46443 27421
rect 46750 27412 46756 27424
rect 46808 27412 46814 27464
rect 47688 27461 47716 27492
rect 48038 27480 48044 27492
rect 48096 27480 48102 27532
rect 47673 27455 47731 27461
rect 47673 27421 47685 27455
rect 47719 27421 47731 27455
rect 47673 27415 47731 27421
rect 47854 27412 47860 27464
rect 47912 27452 47918 27464
rect 48130 27452 48136 27464
rect 47912 27424 48136 27452
rect 47912 27412 47918 27424
rect 48130 27412 48136 27424
rect 48188 27412 48194 27464
rect 48317 27455 48375 27461
rect 48317 27421 48329 27455
rect 48363 27452 48375 27455
rect 48424 27452 48452 27628
rect 49878 27616 49884 27628
rect 49936 27656 49942 27668
rect 50430 27656 50436 27668
rect 49936 27628 50436 27656
rect 49936 27616 49942 27628
rect 50430 27616 50436 27628
rect 50488 27616 50494 27668
rect 51169 27659 51227 27665
rect 51169 27625 51181 27659
rect 51215 27656 51227 27659
rect 51350 27656 51356 27668
rect 51215 27628 51356 27656
rect 51215 27625 51227 27628
rect 51169 27619 51227 27625
rect 51350 27616 51356 27628
rect 51408 27616 51414 27668
rect 51534 27616 51540 27668
rect 51592 27656 51598 27668
rect 52365 27659 52423 27665
rect 52365 27656 52377 27659
rect 51592 27628 52377 27656
rect 51592 27616 51598 27628
rect 52365 27625 52377 27628
rect 52411 27625 52423 27659
rect 52365 27619 52423 27625
rect 53098 27616 53104 27668
rect 53156 27656 53162 27668
rect 58066 27656 58072 27668
rect 53156 27628 58072 27656
rect 53156 27616 53162 27628
rect 58066 27616 58072 27628
rect 58124 27616 58130 27668
rect 48685 27591 48743 27597
rect 48685 27557 48697 27591
rect 48731 27588 48743 27591
rect 48866 27588 48872 27600
rect 48731 27560 48872 27588
rect 48731 27557 48743 27560
rect 48685 27551 48743 27557
rect 48866 27548 48872 27560
rect 48924 27548 48930 27600
rect 49602 27548 49608 27600
rect 49660 27588 49666 27600
rect 50709 27591 50767 27597
rect 50709 27588 50721 27591
rect 49660 27560 50721 27588
rect 49660 27548 49666 27560
rect 50709 27557 50721 27560
rect 50755 27588 50767 27591
rect 53006 27588 53012 27600
rect 50755 27560 52684 27588
rect 52967 27560 53012 27588
rect 50755 27557 50767 27560
rect 50709 27551 50767 27557
rect 48363 27424 48452 27452
rect 48884 27452 48912 27548
rect 49510 27520 49516 27532
rect 49436 27492 49516 27520
rect 49436 27461 49464 27492
rect 49510 27480 49516 27492
rect 49568 27480 49574 27532
rect 51902 27520 51908 27532
rect 51863 27492 51908 27520
rect 51902 27480 51908 27492
rect 51960 27480 51966 27532
rect 49145 27455 49203 27461
rect 49145 27452 49157 27455
rect 48884 27424 49157 27452
rect 48363 27421 48375 27424
rect 48317 27415 48375 27421
rect 49145 27421 49157 27424
rect 49191 27421 49203 27455
rect 49145 27415 49203 27421
rect 49421 27455 49479 27461
rect 49421 27421 49433 27455
rect 49467 27421 49479 27455
rect 49421 27415 49479 27421
rect 49602 27412 49608 27464
rect 49660 27452 49666 27464
rect 50341 27455 50399 27461
rect 50341 27452 50353 27455
rect 49660 27424 50353 27452
rect 49660 27412 49666 27424
rect 50341 27421 50353 27424
rect 50387 27421 50399 27455
rect 50341 27415 50399 27421
rect 50430 27412 50436 27464
rect 50488 27452 50494 27464
rect 50525 27455 50583 27461
rect 50525 27452 50537 27455
rect 50488 27424 50537 27452
rect 50488 27412 50494 27424
rect 50525 27421 50537 27424
rect 50571 27421 50583 27455
rect 50525 27415 50583 27421
rect 50614 27412 50620 27464
rect 50672 27452 50678 27464
rect 51445 27455 51503 27461
rect 51445 27452 51457 27455
rect 50672 27424 51457 27452
rect 50672 27412 50678 27424
rect 51445 27421 51457 27424
rect 51491 27421 51503 27455
rect 51626 27452 51632 27464
rect 51587 27424 51632 27452
rect 51445 27415 51503 27421
rect 51626 27412 51632 27424
rect 51684 27412 51690 27464
rect 52656 27461 52684 27560
rect 53006 27548 53012 27560
rect 53064 27548 53070 27600
rect 57790 27588 57796 27600
rect 57440 27560 57796 27588
rect 53098 27520 53104 27532
rect 53059 27492 53104 27520
rect 53098 27480 53104 27492
rect 53156 27480 53162 27532
rect 53466 27480 53472 27532
rect 53524 27520 53530 27532
rect 57440 27529 57468 27560
rect 57790 27548 57796 27560
rect 57848 27548 57854 27600
rect 54113 27523 54171 27529
rect 54113 27520 54125 27523
rect 53524 27492 54125 27520
rect 53524 27480 53530 27492
rect 54113 27489 54125 27492
rect 54159 27489 54171 27523
rect 57241 27523 57299 27529
rect 57241 27520 57253 27523
rect 54113 27483 54171 27489
rect 55048 27492 57253 27520
rect 51813 27455 51871 27461
rect 51813 27421 51825 27455
rect 51859 27452 51871 27455
rect 52641 27455 52699 27461
rect 51859 27424 52592 27452
rect 51859 27421 51871 27424
rect 51813 27415 51871 27421
rect 34379 27356 35756 27384
rect 34379 27353 34391 27356
rect 34333 27347 34391 27353
rect 36630 27344 36636 27396
rect 36688 27384 36694 27396
rect 39206 27384 39212 27396
rect 36688 27356 38700 27384
rect 39167 27356 39212 27384
rect 36688 27344 36694 27356
rect 33410 27276 33416 27328
rect 33468 27316 33474 27328
rect 33597 27319 33655 27325
rect 33597 27316 33609 27319
rect 33468 27288 33609 27316
rect 33468 27276 33474 27288
rect 33597 27285 33609 27288
rect 33643 27285 33655 27319
rect 33597 27279 33655 27285
rect 38470 27276 38476 27328
rect 38528 27316 38534 27328
rect 38565 27319 38623 27325
rect 38565 27316 38577 27319
rect 38528 27288 38577 27316
rect 38528 27276 38534 27288
rect 38565 27285 38577 27288
rect 38611 27285 38623 27319
rect 38672 27316 38700 27356
rect 39206 27344 39212 27356
rect 39264 27344 39270 27396
rect 42242 27384 42248 27396
rect 39316 27356 42248 27384
rect 39316 27316 39344 27356
rect 42242 27344 42248 27356
rect 42300 27344 42306 27396
rect 42978 27344 42984 27396
rect 43036 27344 43042 27396
rect 44545 27387 44603 27393
rect 44545 27384 44557 27387
rect 43272 27356 44557 27384
rect 38672 27288 39344 27316
rect 38565 27279 38623 27285
rect 41506 27276 41512 27328
rect 41564 27316 41570 27328
rect 43272 27316 43300 27356
rect 44545 27353 44557 27356
rect 44591 27353 44603 27387
rect 44545 27347 44603 27353
rect 45557 27387 45615 27393
rect 45557 27353 45569 27387
rect 45603 27353 45615 27387
rect 45557 27347 45615 27353
rect 46201 27387 46259 27393
rect 46201 27353 46213 27387
rect 46247 27384 46259 27387
rect 47946 27384 47952 27396
rect 46247 27356 47952 27384
rect 46247 27353 46259 27356
rect 46201 27347 46259 27353
rect 43898 27316 43904 27328
rect 41564 27288 43300 27316
rect 43859 27288 43904 27316
rect 41564 27276 41570 27288
rect 43898 27276 43904 27288
rect 43956 27276 43962 27328
rect 44818 27276 44824 27328
rect 44876 27316 44882 27328
rect 45189 27319 45247 27325
rect 45189 27316 45201 27319
rect 44876 27288 45201 27316
rect 44876 27276 44882 27288
rect 45189 27285 45201 27288
rect 45235 27285 45247 27319
rect 45572 27316 45600 27347
rect 47946 27344 47952 27356
rect 48004 27344 48010 27396
rect 48501 27387 48559 27393
rect 48501 27353 48513 27387
rect 48547 27353 48559 27387
rect 48501 27347 48559 27353
rect 47302 27316 47308 27328
rect 45572 27288 47308 27316
rect 45189 27279 45247 27285
rect 47302 27276 47308 27288
rect 47360 27276 47366 27328
rect 47486 27276 47492 27328
rect 47544 27316 47550 27328
rect 48516 27316 48544 27347
rect 48590 27344 48596 27396
rect 48648 27384 48654 27396
rect 49513 27387 49571 27393
rect 49513 27384 49525 27387
rect 48648 27356 49525 27384
rect 48648 27344 48654 27356
rect 49513 27353 49525 27356
rect 49559 27384 49571 27387
rect 51258 27384 51264 27396
rect 49559 27356 51264 27384
rect 49559 27353 49571 27356
rect 49513 27347 49571 27353
rect 51258 27344 51264 27356
rect 51316 27344 51322 27396
rect 49786 27316 49792 27328
rect 47544 27288 49792 27316
rect 47544 27276 47550 27288
rect 49786 27276 49792 27288
rect 49844 27276 49850 27328
rect 50890 27276 50896 27328
rect 50948 27316 50954 27328
rect 51537 27319 51595 27325
rect 51537 27316 51549 27319
rect 50948 27288 51549 27316
rect 50948 27276 50954 27288
rect 51537 27285 51549 27288
rect 51583 27316 51595 27319
rect 52362 27316 52368 27328
rect 51583 27288 52368 27316
rect 51583 27285 51595 27288
rect 51537 27279 51595 27285
rect 52362 27276 52368 27288
rect 52420 27276 52426 27328
rect 52564 27316 52592 27424
rect 52641 27421 52653 27455
rect 52687 27421 52699 27455
rect 52641 27415 52699 27421
rect 52730 27412 52736 27464
rect 52788 27452 52794 27464
rect 53926 27452 53932 27464
rect 52788 27424 52833 27452
rect 53887 27424 53932 27452
rect 52788 27412 52794 27424
rect 53926 27412 53932 27424
rect 53984 27412 53990 27464
rect 54294 27412 54300 27464
rect 54352 27452 54358 27464
rect 54757 27455 54815 27461
rect 54757 27452 54769 27455
rect 54352 27424 54769 27452
rect 54352 27412 54358 27424
rect 54757 27421 54769 27424
rect 54803 27421 54815 27455
rect 54757 27415 54815 27421
rect 54846 27412 54852 27464
rect 54904 27452 54910 27464
rect 54941 27455 54999 27461
rect 54941 27452 54953 27455
rect 54904 27424 54953 27452
rect 54904 27412 54910 27424
rect 54941 27421 54953 27424
rect 54987 27421 54999 27455
rect 54941 27415 54999 27421
rect 52825 27387 52883 27393
rect 52825 27353 52837 27387
rect 52871 27384 52883 27387
rect 55048 27384 55076 27492
rect 57241 27489 57253 27492
rect 57287 27489 57299 27523
rect 57241 27483 57299 27489
rect 57425 27523 57483 27529
rect 57425 27489 57437 27523
rect 57471 27489 57483 27523
rect 57698 27520 57704 27532
rect 57659 27492 57704 27520
rect 57425 27483 57483 27489
rect 57698 27480 57704 27492
rect 57756 27480 57762 27532
rect 55858 27452 55864 27464
rect 55819 27424 55864 27452
rect 55858 27412 55864 27424
rect 55916 27412 55922 27464
rect 56413 27455 56471 27461
rect 56413 27421 56425 27455
rect 56459 27452 56471 27455
rect 56502 27452 56508 27464
rect 56459 27424 56508 27452
rect 56459 27421 56471 27424
rect 56413 27415 56471 27421
rect 56502 27412 56508 27424
rect 56560 27412 56566 27464
rect 57517 27455 57575 27461
rect 57517 27421 57529 27455
rect 57563 27421 57575 27455
rect 57517 27415 57575 27421
rect 57609 27455 57667 27461
rect 57609 27421 57621 27455
rect 57655 27452 57667 27455
rect 58066 27452 58072 27464
rect 57655 27424 58072 27452
rect 57655 27421 57667 27424
rect 57609 27415 57667 27421
rect 52871 27356 55076 27384
rect 55677 27387 55735 27393
rect 52871 27353 52883 27356
rect 52825 27347 52883 27353
rect 55677 27353 55689 27387
rect 55723 27384 55735 27387
rect 56870 27384 56876 27396
rect 55723 27356 56876 27384
rect 55723 27353 55735 27356
rect 55677 27347 55735 27353
rect 56870 27344 56876 27356
rect 56928 27344 56934 27396
rect 57532 27384 57560 27415
rect 58066 27412 58072 27424
rect 58124 27452 58130 27464
rect 58342 27452 58348 27464
rect 58124 27424 58348 27452
rect 58124 27412 58130 27424
rect 58342 27412 58348 27424
rect 58400 27412 58406 27464
rect 58158 27384 58164 27396
rect 57532 27356 58164 27384
rect 58158 27344 58164 27356
rect 58216 27344 58222 27396
rect 53561 27319 53619 27325
rect 53561 27316 53573 27319
rect 52564 27288 53573 27316
rect 53561 27285 53573 27288
rect 53607 27285 53619 27319
rect 53561 27279 53619 27285
rect 54021 27319 54079 27325
rect 54021 27285 54033 27319
rect 54067 27316 54079 27319
rect 54754 27316 54760 27328
rect 54067 27288 54760 27316
rect 54067 27285 54079 27288
rect 54021 27279 54079 27285
rect 54754 27276 54760 27288
rect 54812 27276 54818 27328
rect 54941 27319 54999 27325
rect 54941 27285 54953 27319
rect 54987 27316 54999 27319
rect 55030 27316 55036 27328
rect 54987 27288 55036 27316
rect 54987 27285 54999 27288
rect 54941 27279 54999 27285
rect 55030 27276 55036 27288
rect 55088 27276 55094 27328
rect 55122 27276 55128 27328
rect 55180 27316 55186 27328
rect 55493 27319 55551 27325
rect 55493 27316 55505 27319
rect 55180 27288 55505 27316
rect 55180 27276 55186 27288
rect 55493 27285 55505 27288
rect 55539 27285 55551 27319
rect 58250 27316 58256 27328
rect 58211 27288 58256 27316
rect 55493 27279 55551 27285
rect 58250 27276 58256 27288
rect 58308 27276 58314 27328
rect 1104 27226 58880 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 58880 27226
rect 1104 27152 58880 27174
rect 33778 27072 33784 27124
rect 33836 27112 33842 27124
rect 35621 27115 35679 27121
rect 35621 27112 35633 27115
rect 33836 27084 35633 27112
rect 33836 27072 33842 27084
rect 35621 27081 35633 27084
rect 35667 27081 35679 27115
rect 37461 27115 37519 27121
rect 37461 27112 37473 27115
rect 35621 27075 35679 27081
rect 35728 27084 37473 27112
rect 33410 27044 33416 27056
rect 33371 27016 33416 27044
rect 33410 27004 33416 27016
rect 33468 27004 33474 27056
rect 34146 27004 34152 27056
rect 34204 27004 34210 27056
rect 35342 27004 35348 27056
rect 35400 27044 35406 27056
rect 35728 27044 35756 27084
rect 37461 27081 37473 27084
rect 37507 27081 37519 27115
rect 39022 27112 39028 27124
rect 38983 27084 39028 27112
rect 37461 27075 37519 27081
rect 39022 27072 39028 27084
rect 39080 27072 39086 27124
rect 39577 27115 39635 27121
rect 39577 27081 39589 27115
rect 39623 27112 39635 27115
rect 41322 27112 41328 27124
rect 39623 27084 41328 27112
rect 39623 27081 39635 27084
rect 39577 27075 39635 27081
rect 41322 27072 41328 27084
rect 41380 27072 41386 27124
rect 45554 27112 45560 27124
rect 45515 27084 45560 27112
rect 45554 27072 45560 27084
rect 45612 27072 45618 27124
rect 47857 27115 47915 27121
rect 47857 27081 47869 27115
rect 47903 27112 47915 27115
rect 48038 27112 48044 27124
rect 47903 27084 48044 27112
rect 47903 27081 47915 27084
rect 47857 27075 47915 27081
rect 48038 27072 48044 27084
rect 48096 27072 48102 27124
rect 54297 27115 54355 27121
rect 51046 27084 51764 27112
rect 36817 27047 36875 27053
rect 36817 27044 36829 27047
rect 35400 27016 35756 27044
rect 36004 27016 36829 27044
rect 35400 27004 35406 27016
rect 36004 26988 36032 27016
rect 36817 27013 36829 27016
rect 36863 27013 36875 27047
rect 36817 27007 36875 27013
rect 37182 27004 37188 27056
rect 37240 27044 37246 27056
rect 37921 27047 37979 27053
rect 37240 27016 37780 27044
rect 37240 27004 37246 27016
rect 35986 26976 35992 26988
rect 35947 26948 35992 26976
rect 35986 26936 35992 26948
rect 36044 26936 36050 26988
rect 36081 26979 36139 26985
rect 36081 26945 36093 26979
rect 36127 26976 36139 26979
rect 37752 26976 37780 27016
rect 37921 27013 37933 27047
rect 37967 27044 37979 27047
rect 37967 27016 39528 27044
rect 37967 27013 37979 27016
rect 37921 27007 37979 27013
rect 39500 26988 39528 27016
rect 40770 27004 40776 27056
rect 40828 27004 40834 27056
rect 42518 27004 42524 27056
rect 42576 27044 42582 27056
rect 42797 27047 42855 27053
rect 42797 27044 42809 27047
rect 42576 27016 42809 27044
rect 42576 27004 42582 27016
rect 42797 27013 42809 27016
rect 42843 27013 42855 27047
rect 42797 27007 42855 27013
rect 43901 27047 43959 27053
rect 43901 27013 43913 27047
rect 43947 27044 43959 27047
rect 43990 27044 43996 27056
rect 43947 27016 43996 27044
rect 43947 27013 43959 27016
rect 43901 27007 43959 27013
rect 43990 27004 43996 27016
rect 44048 27004 44054 27056
rect 45094 27044 45100 27056
rect 44560 27016 45100 27044
rect 38470 26976 38476 26988
rect 36127 26948 37688 26976
rect 37752 26948 38476 26976
rect 36127 26945 36139 26948
rect 36081 26939 36139 26945
rect 33137 26911 33195 26917
rect 33137 26877 33149 26911
rect 33183 26908 33195 26911
rect 35161 26911 35219 26917
rect 33183 26880 33272 26908
rect 33183 26877 33195 26880
rect 33137 26871 33195 26877
rect 32858 26732 32864 26784
rect 32916 26772 32922 26784
rect 33244 26772 33272 26880
rect 35161 26877 35173 26911
rect 35207 26908 35219 26911
rect 36096 26908 36124 26939
rect 36262 26908 36268 26920
rect 35207 26880 36124 26908
rect 36223 26880 36268 26908
rect 35207 26877 35219 26880
rect 35161 26871 35219 26877
rect 36262 26868 36268 26880
rect 36320 26868 36326 26920
rect 37550 26840 37556 26852
rect 37511 26812 37556 26840
rect 37550 26800 37556 26812
rect 37608 26800 37614 26852
rect 37660 26840 37688 26948
rect 38470 26936 38476 26948
rect 38528 26936 38534 26988
rect 39482 26976 39488 26988
rect 39395 26948 39488 26976
rect 39482 26936 39488 26948
rect 39540 26936 39546 26988
rect 39669 26979 39727 26985
rect 39669 26945 39681 26979
rect 39715 26976 39727 26979
rect 39942 26976 39948 26988
rect 39715 26948 39948 26976
rect 39715 26945 39727 26948
rect 39669 26939 39727 26945
rect 39942 26936 39948 26948
rect 40000 26936 40006 26988
rect 40678 26976 40684 26988
rect 40639 26948 40684 26976
rect 40678 26936 40684 26948
rect 40736 26936 40742 26988
rect 41138 26976 41144 26988
rect 41099 26948 41144 26976
rect 41138 26936 41144 26948
rect 41196 26936 41202 26988
rect 42978 26936 42984 26988
rect 43036 26976 43042 26988
rect 43073 26979 43131 26985
rect 43073 26976 43085 26979
rect 43036 26948 43085 26976
rect 43036 26936 43042 26948
rect 43073 26945 43085 26948
rect 43119 26976 43131 26979
rect 43625 26979 43683 26985
rect 43625 26976 43637 26979
rect 43119 26948 43637 26976
rect 43119 26945 43131 26948
rect 43073 26939 43131 26945
rect 43625 26945 43637 26948
rect 43671 26945 43683 26979
rect 44450 26976 44456 26988
rect 43625 26939 43683 26945
rect 43732 26948 44456 26976
rect 37734 26868 37740 26920
rect 37792 26908 37798 26920
rect 38194 26908 38200 26920
rect 37792 26880 38200 26908
rect 37792 26868 37798 26880
rect 38194 26868 38200 26880
rect 38252 26908 38258 26920
rect 38749 26911 38807 26917
rect 38749 26908 38761 26911
rect 38252 26880 38761 26908
rect 38252 26868 38258 26880
rect 38749 26877 38761 26880
rect 38795 26908 38807 26911
rect 40218 26908 40224 26920
rect 38795 26880 40224 26908
rect 38795 26877 38807 26880
rect 38749 26871 38807 26877
rect 40218 26868 40224 26880
rect 40276 26868 40282 26920
rect 42426 26868 42432 26920
rect 42484 26908 42490 26920
rect 43732 26908 43760 26948
rect 44450 26936 44456 26948
rect 44508 26936 44514 26988
rect 44560 26985 44588 27016
rect 45094 27004 45100 27016
rect 45152 27004 45158 27056
rect 45646 27004 45652 27056
rect 45704 27044 45710 27056
rect 45704 27016 46428 27044
rect 45704 27004 45710 27016
rect 44545 26979 44603 26985
rect 44545 26945 44557 26979
rect 44591 26945 44603 26979
rect 44545 26939 44603 26945
rect 44637 26979 44695 26985
rect 44637 26945 44649 26979
rect 44683 26945 44695 26979
rect 44818 26976 44824 26988
rect 44779 26948 44824 26976
rect 44637 26939 44695 26945
rect 42484 26880 43760 26908
rect 44652 26908 44680 26939
rect 44818 26936 44824 26948
rect 44876 26936 44882 26988
rect 45738 26936 45744 26988
rect 45796 26976 45802 26988
rect 46201 26979 46259 26985
rect 46201 26976 46213 26979
rect 45796 26948 46213 26976
rect 45796 26936 45802 26948
rect 46201 26945 46213 26948
rect 46247 26976 46259 26979
rect 46290 26976 46296 26988
rect 46247 26948 46296 26976
rect 46247 26945 46259 26948
rect 46201 26939 46259 26945
rect 46290 26936 46296 26948
rect 46348 26936 46354 26988
rect 46400 26985 46428 27016
rect 46658 27004 46664 27056
rect 46716 27044 46722 27056
rect 51046 27044 51074 27084
rect 46716 27016 51074 27044
rect 46716 27004 46722 27016
rect 51258 27004 51264 27056
rect 51316 27044 51322 27056
rect 51316 27016 51580 27044
rect 51316 27004 51322 27016
rect 46385 26979 46443 26985
rect 46385 26945 46397 26979
rect 46431 26976 46443 26979
rect 46842 26976 46848 26988
rect 46431 26948 46848 26976
rect 46431 26945 46443 26948
rect 46385 26939 46443 26945
rect 46842 26936 46848 26948
rect 46900 26976 46906 26988
rect 47029 26979 47087 26985
rect 47029 26976 47041 26979
rect 46900 26948 47041 26976
rect 46900 26936 46906 26948
rect 47029 26945 47041 26948
rect 47075 26945 47087 26979
rect 47029 26939 47087 26945
rect 47213 26979 47271 26985
rect 47213 26945 47225 26979
rect 47259 26945 47271 26979
rect 47213 26939 47271 26945
rect 45756 26908 45784 26936
rect 44652 26880 45784 26908
rect 42484 26868 42490 26880
rect 45830 26868 45836 26920
rect 45888 26908 45894 26920
rect 46750 26908 46756 26920
rect 45888 26880 46756 26908
rect 45888 26868 45894 26880
rect 46750 26868 46756 26880
rect 46808 26908 46814 26920
rect 47228 26908 47256 26939
rect 47670 26936 47676 26988
rect 47728 26976 47734 26988
rect 47765 26979 47823 26985
rect 47765 26976 47777 26979
rect 47728 26948 47777 26976
rect 47728 26936 47734 26948
rect 47765 26945 47777 26948
rect 47811 26945 47823 26979
rect 47765 26939 47823 26945
rect 47949 26979 48007 26985
rect 47949 26945 47961 26979
rect 47995 26945 48007 26979
rect 47949 26939 48007 26945
rect 46808 26880 47256 26908
rect 47964 26908 47992 26939
rect 48130 26936 48136 26988
rect 48188 26976 48194 26988
rect 48777 26979 48835 26985
rect 48777 26976 48789 26979
rect 48188 26948 48789 26976
rect 48188 26936 48194 26948
rect 48777 26945 48789 26948
rect 48823 26945 48835 26979
rect 48777 26939 48835 26945
rect 48958 26936 48964 26988
rect 49016 26976 49022 26988
rect 50062 26976 50068 26988
rect 49016 26948 49061 26976
rect 50023 26948 50068 26976
rect 49016 26936 49022 26948
rect 50062 26936 50068 26948
rect 50120 26936 50126 26988
rect 50154 26936 50160 26988
rect 50212 26976 50218 26988
rect 50338 26976 50344 26988
rect 50212 26948 50257 26976
rect 50299 26948 50344 26976
rect 50212 26936 50218 26948
rect 50338 26936 50344 26948
rect 50396 26936 50402 26988
rect 50433 26979 50491 26985
rect 50433 26945 50445 26979
rect 50479 26945 50491 26979
rect 50433 26939 50491 26945
rect 48866 26908 48872 26920
rect 47964 26880 48872 26908
rect 46808 26868 46814 26880
rect 48866 26868 48872 26880
rect 48924 26868 48930 26920
rect 49050 26868 49056 26920
rect 49108 26908 49114 26920
rect 50448 26908 50476 26939
rect 50522 26936 50528 26988
rect 50580 26976 50586 26988
rect 50580 26948 50625 26976
rect 50580 26936 50586 26948
rect 51166 26936 51172 26988
rect 51224 26976 51230 26988
rect 51353 26979 51411 26985
rect 51353 26976 51365 26979
rect 51224 26948 51365 26976
rect 51224 26936 51230 26948
rect 51353 26945 51365 26948
rect 51399 26945 51411 26979
rect 51353 26939 51411 26945
rect 51445 26979 51503 26985
rect 51445 26945 51457 26979
rect 51491 26945 51503 26979
rect 51445 26939 51503 26945
rect 50890 26908 50896 26920
rect 49108 26880 50896 26908
rect 49108 26868 49114 26880
rect 50890 26868 50896 26880
rect 50948 26868 50954 26920
rect 51460 26908 51488 26939
rect 51046 26880 51488 26908
rect 51552 26908 51580 27016
rect 51736 26985 51764 27084
rect 54297 27081 54309 27115
rect 54343 27112 54355 27115
rect 54478 27112 54484 27124
rect 54343 27084 54484 27112
rect 54343 27081 54355 27084
rect 54297 27075 54355 27081
rect 54478 27072 54484 27084
rect 54536 27072 54542 27124
rect 54754 27112 54760 27124
rect 54715 27084 54760 27112
rect 54754 27072 54760 27084
rect 54812 27072 54818 27124
rect 55953 27115 56011 27121
rect 54864 27084 55812 27112
rect 53190 27044 53196 27056
rect 52472 27016 53196 27044
rect 51721 26979 51779 26985
rect 51721 26945 51733 26979
rect 51767 26976 51779 26979
rect 52362 26976 52368 26988
rect 51767 26948 52368 26976
rect 51767 26945 51779 26948
rect 51721 26939 51779 26945
rect 52362 26936 52368 26948
rect 52420 26936 52426 26988
rect 52472 26908 52500 27016
rect 53190 27004 53196 27016
rect 53248 27044 53254 27056
rect 54864 27044 54892 27084
rect 55030 27044 55036 27056
rect 53248 27016 54892 27044
rect 54991 27016 55036 27044
rect 53248 27004 53254 27016
rect 55030 27004 55036 27016
rect 55088 27004 55094 27056
rect 55122 27004 55128 27056
rect 55180 27044 55186 27056
rect 55784 27053 55812 27084
rect 55953 27081 55965 27115
rect 55999 27112 56011 27115
rect 56870 27112 56876 27124
rect 55999 27084 56876 27112
rect 55999 27081 56011 27084
rect 55953 27075 56011 27081
rect 56870 27072 56876 27084
rect 56928 27072 56934 27124
rect 55769 27047 55827 27053
rect 55180 27016 55225 27044
rect 55180 27004 55186 27016
rect 55769 27013 55781 27047
rect 55815 27013 55827 27047
rect 55769 27007 55827 27013
rect 55858 27004 55864 27056
rect 55916 27044 55922 27056
rect 56597 27047 56655 27053
rect 55916 27016 56088 27044
rect 55916 27004 55922 27016
rect 53377 26979 53435 26985
rect 53377 26945 53389 26979
rect 53423 26976 53435 26979
rect 53558 26976 53564 26988
rect 53423 26948 53564 26976
rect 53423 26945 53435 26948
rect 53377 26939 53435 26945
rect 53558 26936 53564 26948
rect 53616 26936 53622 26988
rect 54662 26936 54668 26988
rect 54720 26976 54726 26988
rect 56060 26985 56088 27016
rect 56597 27013 56609 27047
rect 56643 27044 56655 27047
rect 56686 27044 56692 27056
rect 56643 27016 56692 27044
rect 56643 27013 56655 27016
rect 56597 27007 56655 27013
rect 56686 27004 56692 27016
rect 56744 27044 56750 27056
rect 57882 27044 57888 27056
rect 56744 27016 57888 27044
rect 56744 27004 56750 27016
rect 57882 27004 57888 27016
rect 57940 27004 57946 27056
rect 54941 26979 54999 26985
rect 54941 26976 54953 26979
rect 54720 26948 54953 26976
rect 54720 26936 54726 26948
rect 54941 26945 54953 26948
rect 54987 26945 54999 26979
rect 54941 26939 54999 26945
rect 55309 26979 55367 26985
rect 55309 26945 55321 26979
rect 55355 26945 55367 26979
rect 55309 26939 55367 26945
rect 56045 26979 56103 26985
rect 56045 26945 56057 26979
rect 56091 26945 56103 26979
rect 56045 26939 56103 26945
rect 53282 26908 53288 26920
rect 51552 26880 52500 26908
rect 53243 26880 53288 26908
rect 37660 26812 41414 26840
rect 34606 26772 34612 26784
rect 32916 26744 34612 26772
rect 32916 26732 32922 26744
rect 34606 26732 34612 26744
rect 34664 26732 34670 26784
rect 38562 26772 38568 26784
rect 38523 26744 38568 26772
rect 38562 26732 38568 26744
rect 38620 26732 38626 26784
rect 41386 26772 41414 26812
rect 46382 26800 46388 26852
rect 46440 26840 46446 26852
rect 46477 26843 46535 26849
rect 46477 26840 46489 26843
rect 46440 26812 46489 26840
rect 46440 26800 46446 26812
rect 46477 26809 46489 26812
rect 46523 26840 46535 26843
rect 46566 26840 46572 26852
rect 46523 26812 46572 26840
rect 46523 26809 46535 26812
rect 46477 26803 46535 26809
rect 46566 26800 46572 26812
rect 46624 26800 46630 26852
rect 50709 26843 50767 26849
rect 50709 26809 50721 26843
rect 50755 26840 50767 26843
rect 51046 26840 51074 26880
rect 53282 26868 53288 26880
rect 53340 26868 53346 26920
rect 55324 26908 55352 26939
rect 55324 26880 55812 26908
rect 50755 26812 51074 26840
rect 53745 26843 53803 26849
rect 50755 26809 50767 26812
rect 50709 26803 50767 26809
rect 53745 26809 53757 26843
rect 53791 26840 53803 26843
rect 54294 26840 54300 26852
rect 53791 26812 54300 26840
rect 53791 26809 53803 26812
rect 53745 26803 53803 26809
rect 54294 26800 54300 26812
rect 54352 26800 54358 26852
rect 55784 26849 55812 26880
rect 55769 26843 55827 26849
rect 55769 26809 55781 26843
rect 55815 26809 55827 26843
rect 55769 26803 55827 26809
rect 43622 26772 43628 26784
rect 41386 26744 43628 26772
rect 43622 26732 43628 26744
rect 43680 26732 43686 26784
rect 45005 26775 45063 26781
rect 45005 26741 45017 26775
rect 45051 26772 45063 26775
rect 47026 26772 47032 26784
rect 45051 26744 47032 26772
rect 45051 26741 45063 26744
rect 45005 26735 45063 26741
rect 47026 26732 47032 26744
rect 47084 26732 47090 26784
rect 47121 26775 47179 26781
rect 47121 26741 47133 26775
rect 47167 26772 47179 26775
rect 48130 26772 48136 26784
rect 47167 26744 48136 26772
rect 47167 26741 47179 26744
rect 47121 26735 47179 26741
rect 48130 26732 48136 26744
rect 48188 26732 48194 26784
rect 49145 26775 49203 26781
rect 49145 26741 49157 26775
rect 49191 26772 49203 26775
rect 49602 26772 49608 26784
rect 49191 26744 49608 26772
rect 49191 26741 49203 26744
rect 49145 26735 49203 26741
rect 49602 26732 49608 26744
rect 49660 26732 49666 26784
rect 51169 26775 51227 26781
rect 51169 26741 51181 26775
rect 51215 26772 51227 26775
rect 51258 26772 51264 26784
rect 51215 26744 51264 26772
rect 51215 26741 51227 26744
rect 51169 26735 51227 26741
rect 51258 26732 51264 26744
rect 51316 26732 51322 26784
rect 51626 26772 51632 26784
rect 51587 26744 51632 26772
rect 51626 26732 51632 26744
rect 51684 26732 51690 26784
rect 52178 26772 52184 26784
rect 52139 26744 52184 26772
rect 52178 26732 52184 26744
rect 52236 26772 52242 26784
rect 53466 26772 53472 26784
rect 52236 26744 53472 26772
rect 52236 26732 52242 26744
rect 53466 26732 53472 26744
rect 53524 26732 53530 26784
rect 53558 26732 53564 26784
rect 53616 26772 53622 26784
rect 56594 26772 56600 26784
rect 53616 26744 56600 26772
rect 53616 26732 53622 26744
rect 56594 26732 56600 26744
rect 56652 26772 56658 26784
rect 57149 26775 57207 26781
rect 57149 26772 57161 26775
rect 56652 26744 57161 26772
rect 56652 26732 56658 26744
rect 57149 26741 57161 26744
rect 57195 26741 57207 26775
rect 58066 26772 58072 26784
rect 58027 26744 58072 26772
rect 57149 26735 57207 26741
rect 58066 26732 58072 26744
rect 58124 26732 58130 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 2406 26528 2412 26580
rect 2464 26568 2470 26580
rect 31665 26571 31723 26577
rect 2464 26540 26234 26568
rect 2464 26528 2470 26540
rect 26206 26500 26234 26540
rect 31665 26537 31677 26571
rect 31711 26568 31723 26571
rect 32306 26568 32312 26580
rect 31711 26540 32312 26568
rect 31711 26537 31723 26540
rect 31665 26531 31723 26537
rect 32306 26528 32312 26540
rect 32364 26568 32370 26580
rect 32858 26568 32864 26580
rect 32364 26540 32864 26568
rect 32364 26528 32370 26540
rect 32858 26528 32864 26540
rect 32916 26528 32922 26580
rect 34146 26528 34152 26580
rect 34204 26568 34210 26580
rect 34241 26571 34299 26577
rect 34241 26568 34253 26571
rect 34204 26540 34253 26568
rect 34204 26528 34210 26540
rect 34241 26537 34253 26540
rect 34287 26537 34299 26571
rect 36630 26568 36636 26580
rect 36591 26540 36636 26568
rect 34241 26531 34299 26537
rect 36630 26528 36636 26540
rect 36688 26528 36694 26580
rect 37921 26571 37979 26577
rect 37921 26537 37933 26571
rect 37967 26568 37979 26571
rect 38930 26568 38936 26580
rect 37967 26540 38936 26568
rect 37967 26537 37979 26540
rect 37921 26531 37979 26537
rect 38930 26528 38936 26540
rect 38988 26528 38994 26580
rect 39482 26528 39488 26580
rect 39540 26568 39546 26580
rect 40037 26571 40095 26577
rect 40037 26568 40049 26571
rect 39540 26540 40049 26568
rect 39540 26528 39546 26540
rect 40037 26537 40049 26540
rect 40083 26537 40095 26571
rect 40037 26531 40095 26537
rect 40221 26571 40279 26577
rect 40221 26537 40233 26571
rect 40267 26537 40279 26571
rect 40221 26531 40279 26537
rect 41877 26571 41935 26577
rect 41877 26537 41889 26571
rect 41923 26568 41935 26571
rect 44082 26568 44088 26580
rect 41923 26540 44088 26568
rect 41923 26537 41935 26540
rect 41877 26531 41935 26537
rect 40126 26500 40132 26512
rect 26206 26472 35020 26500
rect 34698 26392 34704 26444
rect 34756 26432 34762 26444
rect 34885 26435 34943 26441
rect 34885 26432 34897 26435
rect 34756 26404 34897 26432
rect 34756 26392 34762 26404
rect 34885 26401 34897 26404
rect 34931 26401 34943 26435
rect 34992 26432 35020 26472
rect 36188 26472 40132 26500
rect 36188 26432 36216 26472
rect 40126 26460 40132 26472
rect 40184 26460 40190 26512
rect 40236 26444 40264 26531
rect 44082 26528 44088 26540
rect 44140 26528 44146 26580
rect 45281 26571 45339 26577
rect 45281 26537 45293 26571
rect 45327 26568 45339 26571
rect 45830 26568 45836 26580
rect 45327 26540 45836 26568
rect 45327 26537 45339 26540
rect 45281 26531 45339 26537
rect 45830 26528 45836 26540
rect 45888 26528 45894 26580
rect 46842 26528 46848 26580
rect 46900 26568 46906 26580
rect 47029 26571 47087 26577
rect 47029 26568 47041 26571
rect 46900 26540 47041 26568
rect 46900 26528 46906 26540
rect 47029 26537 47041 26540
rect 47075 26537 47087 26571
rect 50433 26571 50491 26577
rect 47029 26531 47087 26537
rect 47688 26540 49556 26568
rect 47688 26512 47716 26540
rect 42426 26500 42432 26512
rect 42387 26472 42432 26500
rect 42426 26460 42432 26472
rect 42484 26460 42490 26512
rect 47210 26500 47216 26512
rect 45204 26472 47216 26500
rect 34992 26404 36216 26432
rect 34885 26395 34943 26401
rect 36446 26392 36452 26444
rect 36504 26432 36510 26444
rect 37553 26435 37611 26441
rect 37553 26432 37565 26435
rect 36504 26404 37565 26432
rect 36504 26392 36510 26404
rect 37553 26401 37565 26404
rect 37599 26432 37611 26435
rect 38562 26432 38568 26444
rect 37599 26404 38568 26432
rect 37599 26401 37611 26404
rect 37553 26395 37611 26401
rect 38562 26392 38568 26404
rect 38620 26392 38626 26444
rect 39206 26432 39212 26444
rect 39167 26404 39212 26432
rect 39206 26392 39212 26404
rect 39264 26392 39270 26444
rect 40218 26392 40224 26444
rect 40276 26392 40282 26444
rect 40310 26392 40316 26444
rect 40368 26432 40374 26444
rect 41138 26432 41144 26444
rect 40368 26404 41144 26432
rect 40368 26392 40374 26404
rect 41138 26392 41144 26404
rect 41196 26392 41202 26444
rect 41322 26432 41328 26444
rect 41283 26404 41328 26432
rect 41322 26392 41328 26404
rect 41380 26392 41386 26444
rect 32950 26364 32956 26376
rect 32911 26336 32956 26364
rect 32950 26324 32956 26336
rect 33008 26324 33014 26376
rect 34149 26367 34207 26373
rect 34149 26333 34161 26367
rect 34195 26364 34207 26367
rect 34790 26364 34796 26376
rect 34195 26336 34796 26364
rect 34195 26333 34207 26336
rect 34149 26327 34207 26333
rect 34790 26324 34796 26336
rect 34848 26324 34854 26376
rect 37642 26364 37648 26376
rect 37603 26336 37648 26364
rect 37642 26324 37648 26336
rect 37700 26324 37706 26376
rect 37737 26367 37795 26373
rect 37737 26333 37749 26367
rect 37783 26333 37795 26367
rect 37737 26327 37795 26333
rect 39485 26367 39543 26373
rect 39485 26333 39497 26367
rect 39531 26364 39543 26367
rect 39666 26364 39672 26376
rect 39531 26336 39672 26364
rect 39531 26333 39543 26336
rect 39485 26327 39543 26333
rect 35158 26296 35164 26308
rect 35119 26268 35164 26296
rect 35158 26256 35164 26268
rect 35216 26256 35222 26308
rect 36170 26256 36176 26308
rect 36228 26256 36234 26308
rect 36538 26256 36544 26308
rect 36596 26296 36602 26308
rect 37182 26296 37188 26308
rect 36596 26268 37188 26296
rect 36596 26256 36602 26268
rect 37182 26256 37188 26268
rect 37240 26296 37246 26308
rect 37752 26296 37780 26327
rect 39666 26324 39672 26336
rect 39724 26324 39730 26376
rect 40494 26324 40500 26376
rect 40552 26364 40558 26376
rect 40589 26367 40647 26373
rect 40589 26364 40601 26367
rect 40552 26336 40601 26364
rect 40552 26324 40558 26336
rect 40589 26333 40601 26336
rect 40635 26364 40647 26367
rect 40678 26364 40684 26376
rect 40635 26336 40684 26364
rect 40635 26333 40647 26336
rect 40589 26327 40647 26333
rect 40678 26324 40684 26336
rect 40736 26324 40742 26376
rect 41417 26367 41475 26373
rect 41417 26333 41429 26367
rect 41463 26364 41475 26367
rect 41506 26364 41512 26376
rect 41463 26336 41512 26364
rect 41463 26333 41475 26336
rect 41417 26327 41475 26333
rect 41432 26296 41460 26327
rect 41506 26324 41512 26336
rect 41564 26324 41570 26376
rect 42444 26296 42472 26460
rect 42702 26392 42708 26444
rect 42760 26432 42766 26444
rect 44177 26435 44235 26441
rect 44177 26432 44189 26435
rect 42760 26404 44189 26432
rect 42760 26392 42766 26404
rect 44177 26401 44189 26404
rect 44223 26401 44235 26435
rect 44177 26395 44235 26401
rect 45002 26324 45008 26376
rect 45060 26364 45066 26376
rect 45204 26373 45232 26472
rect 47210 26460 47216 26472
rect 47268 26500 47274 26512
rect 47670 26500 47676 26512
rect 47268 26472 47676 26500
rect 47268 26460 47274 26472
rect 47670 26460 47676 26472
rect 47728 26460 47734 26512
rect 47857 26503 47915 26509
rect 47857 26469 47869 26503
rect 47903 26500 47915 26503
rect 48866 26500 48872 26512
rect 47903 26472 48872 26500
rect 47903 26469 47915 26472
rect 47857 26463 47915 26469
rect 48866 26460 48872 26472
rect 48924 26460 48930 26512
rect 46474 26432 46480 26444
rect 46435 26404 46480 26432
rect 46474 26392 46480 26404
rect 46532 26392 46538 26444
rect 46750 26392 46756 26444
rect 46808 26432 46814 26444
rect 48041 26435 48099 26441
rect 46808 26404 47808 26432
rect 46808 26392 46814 26404
rect 45189 26367 45247 26373
rect 45189 26364 45201 26367
rect 45060 26336 45201 26364
rect 45060 26324 45066 26336
rect 45189 26333 45201 26336
rect 45235 26333 45247 26367
rect 45189 26327 45247 26333
rect 47029 26367 47087 26373
rect 47029 26333 47041 26367
rect 47075 26364 47087 26367
rect 47118 26364 47124 26376
rect 47075 26336 47124 26364
rect 47075 26333 47087 26336
rect 47029 26327 47087 26333
rect 47118 26324 47124 26336
rect 47176 26324 47182 26376
rect 47213 26367 47271 26373
rect 47213 26333 47225 26367
rect 47259 26364 47271 26367
rect 47486 26364 47492 26376
rect 47259 26336 47492 26364
rect 47259 26333 47271 26336
rect 47213 26327 47271 26333
rect 43622 26296 43628 26308
rect 37240 26268 37780 26296
rect 37844 26268 41460 26296
rect 41524 26268 42472 26296
rect 43470 26268 43628 26296
rect 37240 26256 37246 26268
rect 35986 26188 35992 26240
rect 36044 26228 36050 26240
rect 37844 26228 37872 26268
rect 36044 26200 37872 26228
rect 36044 26188 36050 26200
rect 38010 26188 38016 26240
rect 38068 26228 38074 26240
rect 40310 26228 40316 26240
rect 38068 26200 40316 26228
rect 38068 26188 38074 26200
rect 40310 26188 40316 26200
rect 40368 26188 40374 26240
rect 41524 26237 41552 26268
rect 43622 26256 43628 26268
rect 43680 26256 43686 26308
rect 43898 26296 43904 26308
rect 43859 26268 43904 26296
rect 43898 26256 43904 26268
rect 43956 26256 43962 26308
rect 45922 26256 45928 26308
rect 45980 26296 45986 26308
rect 46293 26299 46351 26305
rect 46293 26296 46305 26299
rect 45980 26268 46305 26296
rect 45980 26256 45986 26268
rect 46293 26265 46305 26268
rect 46339 26296 46351 26299
rect 47228 26296 47256 26327
rect 47486 26324 47492 26336
rect 47544 26324 47550 26376
rect 47780 26373 47808 26404
rect 48041 26401 48053 26435
rect 48087 26432 48099 26435
rect 48222 26432 48228 26444
rect 48087 26404 48228 26432
rect 48087 26401 48099 26404
rect 48041 26395 48099 26401
rect 48222 26392 48228 26404
rect 48280 26392 48286 26444
rect 49528 26432 49556 26540
rect 50433 26537 50445 26571
rect 50479 26568 50491 26571
rect 50614 26568 50620 26580
rect 50479 26540 50620 26568
rect 50479 26537 50491 26540
rect 50433 26531 50491 26537
rect 50614 26528 50620 26540
rect 50672 26528 50678 26580
rect 52362 26568 52368 26580
rect 52323 26540 52368 26568
rect 52362 26528 52368 26540
rect 52420 26528 52426 26580
rect 52914 26568 52920 26580
rect 52875 26540 52920 26568
rect 52914 26528 52920 26540
rect 52972 26528 52978 26580
rect 53558 26568 53564 26580
rect 53519 26540 53564 26568
rect 53558 26528 53564 26540
rect 53616 26528 53622 26580
rect 54294 26568 54300 26580
rect 54255 26540 54300 26568
rect 54294 26528 54300 26540
rect 54352 26528 54358 26580
rect 54662 26568 54668 26580
rect 54623 26540 54668 26568
rect 54662 26528 54668 26540
rect 54720 26528 54726 26580
rect 55585 26571 55643 26577
rect 55585 26537 55597 26571
rect 55631 26568 55643 26571
rect 56318 26568 56324 26580
rect 55631 26540 56324 26568
rect 55631 26537 55643 26540
rect 55585 26531 55643 26537
rect 56318 26528 56324 26540
rect 56376 26528 56382 26580
rect 56686 26568 56692 26580
rect 56647 26540 56692 26568
rect 56686 26528 56692 26540
rect 56744 26528 56750 26580
rect 54478 26460 54484 26512
rect 54536 26500 54542 26512
rect 56045 26503 56103 26509
rect 56045 26500 56057 26503
rect 54536 26472 56057 26500
rect 54536 26460 54542 26472
rect 56045 26469 56057 26472
rect 56091 26469 56103 26503
rect 56045 26463 56103 26469
rect 49694 26432 49700 26444
rect 49528 26404 49700 26432
rect 47765 26367 47823 26373
rect 47765 26333 47777 26367
rect 47811 26333 47823 26367
rect 47765 26327 47823 26333
rect 48130 26324 48136 26376
rect 48188 26364 48194 26376
rect 48501 26367 48559 26373
rect 48501 26364 48513 26367
rect 48188 26336 48513 26364
rect 48188 26324 48194 26336
rect 48501 26333 48513 26336
rect 48547 26333 48559 26367
rect 48501 26327 48559 26333
rect 48685 26367 48743 26373
rect 48685 26333 48697 26367
rect 48731 26364 48743 26367
rect 48958 26364 48964 26376
rect 48731 26336 48964 26364
rect 48731 26333 48743 26336
rect 48685 26327 48743 26333
rect 46339 26268 47256 26296
rect 46339 26265 46351 26268
rect 46293 26259 46351 26265
rect 47670 26256 47676 26308
rect 47728 26296 47734 26308
rect 48041 26299 48099 26305
rect 48041 26296 48053 26299
rect 47728 26268 48053 26296
rect 47728 26256 47734 26268
rect 48041 26265 48053 26268
rect 48087 26265 48099 26299
rect 48041 26259 48099 26265
rect 48314 26256 48320 26308
rect 48372 26296 48378 26308
rect 48700 26296 48728 26327
rect 48958 26324 48964 26336
rect 49016 26364 49022 26376
rect 49145 26367 49203 26373
rect 49145 26364 49157 26367
rect 49016 26336 49157 26364
rect 49016 26324 49022 26336
rect 49145 26333 49157 26336
rect 49191 26333 49203 26367
rect 49326 26364 49332 26376
rect 49287 26336 49332 26364
rect 49145 26327 49203 26333
rect 49326 26324 49332 26336
rect 49384 26324 49390 26376
rect 49528 26373 49556 26404
rect 49694 26392 49700 26404
rect 49752 26392 49758 26444
rect 54205 26435 54263 26441
rect 54205 26401 54217 26435
rect 54251 26432 54263 26435
rect 54846 26432 54852 26444
rect 54251 26404 54852 26432
rect 54251 26401 54263 26404
rect 54205 26395 54263 26401
rect 54846 26392 54852 26404
rect 54904 26392 54910 26444
rect 49421 26367 49479 26373
rect 49421 26333 49433 26367
rect 49467 26333 49479 26367
rect 49421 26327 49479 26333
rect 49513 26367 49571 26373
rect 49513 26333 49525 26367
rect 49559 26333 49571 26367
rect 49513 26327 49571 26333
rect 48372 26268 48728 26296
rect 48372 26256 48378 26268
rect 48774 26256 48780 26308
rect 48832 26296 48838 26308
rect 49436 26296 49464 26327
rect 49602 26324 49608 26376
rect 49660 26364 49666 26376
rect 50341 26367 50399 26373
rect 50341 26364 50353 26367
rect 49660 26336 50353 26364
rect 49660 26324 49666 26336
rect 50341 26333 50353 26336
rect 50387 26333 50399 26367
rect 50522 26364 50528 26376
rect 50483 26336 50528 26364
rect 50341 26327 50399 26333
rect 50522 26324 50528 26336
rect 50580 26324 50586 26376
rect 50985 26367 51043 26373
rect 50985 26333 50997 26367
rect 51031 26364 51043 26367
rect 51074 26364 51080 26376
rect 51031 26336 51080 26364
rect 51031 26333 51043 26336
rect 50985 26327 51043 26333
rect 51074 26324 51080 26336
rect 51132 26324 51138 26376
rect 51258 26373 51264 26376
rect 51252 26364 51264 26373
rect 51219 26336 51264 26364
rect 51252 26327 51264 26336
rect 51258 26324 51264 26327
rect 51316 26324 51322 26376
rect 52270 26324 52276 26376
rect 52328 26364 52334 26376
rect 54481 26367 54539 26373
rect 54481 26364 54493 26367
rect 52328 26336 54493 26364
rect 52328 26324 52334 26336
rect 54481 26333 54493 26336
rect 54527 26333 54539 26367
rect 54481 26327 54539 26333
rect 48832 26268 49464 26296
rect 49789 26299 49847 26305
rect 48832 26256 48838 26268
rect 49789 26265 49801 26299
rect 49835 26296 49847 26299
rect 51166 26296 51172 26308
rect 49835 26268 51172 26296
rect 49835 26265 49847 26268
rect 49789 26259 49847 26265
rect 51166 26256 51172 26268
rect 51224 26256 51230 26308
rect 57241 26299 57299 26305
rect 57241 26296 57253 26299
rect 52840 26268 53604 26296
rect 41509 26231 41567 26237
rect 41509 26197 41521 26231
rect 41555 26197 41567 26231
rect 45830 26228 45836 26240
rect 45791 26200 45836 26228
rect 41509 26191 41567 26197
rect 45830 26188 45836 26200
rect 45888 26188 45894 26240
rect 46201 26231 46259 26237
rect 46201 26197 46213 26231
rect 46247 26228 46259 26231
rect 46382 26228 46388 26240
rect 46247 26200 46388 26228
rect 46247 26197 46259 26200
rect 46201 26191 46259 26197
rect 46382 26188 46388 26200
rect 46440 26188 46446 26240
rect 48685 26231 48743 26237
rect 48685 26197 48697 26231
rect 48731 26228 48743 26231
rect 50522 26228 50528 26240
rect 48731 26200 50528 26228
rect 48731 26197 48743 26200
rect 48685 26191 48743 26197
rect 50522 26188 50528 26200
rect 50580 26188 50586 26240
rect 50982 26188 50988 26240
rect 51040 26228 51046 26240
rect 52840 26228 52868 26268
rect 51040 26200 52868 26228
rect 53576 26228 53604 26268
rect 55968 26268 57253 26296
rect 55968 26228 55996 26268
rect 57241 26265 57253 26268
rect 57287 26296 57299 26299
rect 58066 26296 58072 26308
rect 57287 26268 58072 26296
rect 57287 26265 57299 26268
rect 57241 26259 57299 26265
rect 58066 26256 58072 26268
rect 58124 26256 58130 26308
rect 53576 26200 55996 26228
rect 51040 26188 51046 26200
rect 1104 26138 58880 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 58880 26138
rect 1104 26064 58880 26086
rect 34517 26027 34575 26033
rect 34517 25993 34529 26027
rect 34563 26024 34575 26027
rect 34698 26024 34704 26036
rect 34563 25996 34704 26024
rect 34563 25993 34575 25996
rect 34517 25987 34575 25993
rect 34698 25984 34704 25996
rect 34756 25984 34762 26036
rect 35158 26024 35164 26036
rect 35119 25996 35164 26024
rect 35158 25984 35164 25996
rect 35216 25984 35222 26036
rect 36262 25984 36268 26036
rect 36320 26024 36326 26036
rect 37461 26027 37519 26033
rect 37461 26024 37473 26027
rect 36320 25996 37473 26024
rect 36320 25984 36326 25996
rect 37461 25993 37473 25996
rect 37507 25993 37519 26027
rect 37461 25987 37519 25993
rect 39114 25984 39120 26036
rect 39172 26024 39178 26036
rect 39577 26027 39635 26033
rect 39577 26024 39589 26027
rect 39172 25996 39589 26024
rect 39172 25984 39178 25996
rect 39577 25993 39589 25996
rect 39623 26024 39635 26027
rect 41414 26024 41420 26036
rect 39623 25996 41420 26024
rect 39623 25993 39635 25996
rect 39577 25987 39635 25993
rect 41414 25984 41420 25996
rect 41472 25984 41478 26036
rect 42242 25984 42248 26036
rect 42300 26024 42306 26036
rect 42610 26024 42616 26036
rect 42300 25996 42616 26024
rect 42300 25984 42306 25996
rect 42610 25984 42616 25996
rect 42668 26024 42674 26036
rect 43622 26024 43628 26036
rect 42668 25996 42932 26024
rect 43583 25996 43628 26024
rect 42668 25984 42674 25996
rect 36173 25959 36231 25965
rect 36173 25925 36185 25959
rect 36219 25956 36231 25959
rect 36630 25956 36636 25968
rect 36219 25928 36636 25956
rect 36219 25925 36231 25928
rect 36173 25919 36231 25925
rect 36630 25916 36636 25928
rect 36688 25916 36694 25968
rect 38010 25956 38016 25968
rect 37660 25928 38016 25956
rect 34977 25891 35035 25897
rect 34977 25857 34989 25891
rect 35023 25888 35035 25891
rect 35023 25860 35848 25888
rect 35023 25857 35035 25860
rect 34977 25851 35035 25857
rect 35820 25761 35848 25860
rect 37458 25848 37464 25900
rect 37516 25888 37522 25900
rect 37660 25897 37688 25928
rect 38010 25916 38016 25928
rect 38068 25916 38074 25968
rect 40129 25959 40187 25965
rect 40129 25956 40141 25959
rect 38396 25928 40141 25956
rect 38396 25897 38424 25928
rect 40129 25925 40141 25928
rect 40175 25956 40187 25959
rect 41230 25956 41236 25968
rect 40175 25928 41236 25956
rect 40175 25925 40187 25928
rect 40129 25919 40187 25925
rect 41230 25916 41236 25928
rect 41288 25916 41294 25968
rect 42904 25965 42932 25996
rect 43622 25984 43628 25996
rect 43680 25984 43686 26036
rect 46290 26024 46296 26036
rect 46251 25996 46296 26024
rect 46290 25984 46296 25996
rect 46348 25984 46354 26036
rect 46934 26024 46940 26036
rect 46895 25996 46940 26024
rect 46934 25984 46940 25996
rect 46992 25984 46998 26036
rect 49510 26024 49516 26036
rect 49068 25996 49516 26024
rect 42889 25959 42947 25965
rect 42889 25925 42901 25959
rect 42935 25925 42947 25959
rect 47118 25956 47124 25968
rect 42889 25919 42947 25925
rect 46124 25928 47124 25956
rect 37645 25891 37703 25897
rect 37645 25888 37657 25891
rect 37516 25860 37657 25888
rect 37516 25848 37522 25860
rect 37645 25857 37657 25860
rect 37691 25857 37703 25891
rect 37645 25851 37703 25857
rect 37921 25891 37979 25897
rect 37921 25857 37933 25891
rect 37967 25888 37979 25891
rect 38381 25891 38439 25897
rect 37967 25860 38332 25888
rect 37967 25857 37979 25860
rect 37921 25851 37979 25857
rect 35986 25820 35992 25832
rect 35912 25792 35992 25820
rect 35805 25755 35863 25761
rect 35805 25721 35817 25755
rect 35851 25721 35863 25755
rect 35805 25715 35863 25721
rect 34790 25644 34796 25696
rect 34848 25684 34854 25696
rect 35912 25684 35940 25792
rect 35986 25780 35992 25792
rect 36044 25820 36050 25832
rect 36265 25823 36323 25829
rect 36265 25820 36277 25823
rect 36044 25792 36277 25820
rect 36044 25780 36050 25792
rect 36265 25789 36277 25792
rect 36311 25789 36323 25823
rect 36265 25783 36323 25789
rect 36449 25823 36507 25829
rect 36449 25789 36461 25823
rect 36495 25789 36507 25823
rect 36449 25783 36507 25789
rect 37829 25823 37887 25829
rect 37829 25789 37841 25823
rect 37875 25820 37887 25823
rect 38010 25820 38016 25832
rect 37875 25792 38016 25820
rect 37875 25789 37887 25792
rect 37829 25783 37887 25789
rect 36464 25752 36492 25783
rect 38010 25780 38016 25792
rect 38068 25780 38074 25832
rect 38304 25820 38332 25860
rect 38381 25857 38393 25891
rect 38427 25857 38439 25891
rect 38381 25851 38439 25857
rect 38565 25891 38623 25897
rect 38565 25857 38577 25891
rect 38611 25857 38623 25891
rect 38565 25851 38623 25857
rect 38304 25792 38516 25820
rect 36464 25724 37964 25752
rect 37936 25693 37964 25724
rect 34848 25656 35940 25684
rect 37921 25687 37979 25693
rect 34848 25644 34854 25656
rect 37921 25653 37933 25687
rect 37967 25684 37979 25687
rect 38102 25684 38108 25696
rect 37967 25656 38108 25684
rect 37967 25653 37979 25656
rect 37921 25647 37979 25653
rect 38102 25644 38108 25656
rect 38160 25644 38166 25696
rect 38488 25693 38516 25792
rect 38580 25752 38608 25851
rect 38654 25848 38660 25900
rect 38712 25888 38718 25900
rect 39301 25891 39359 25897
rect 39301 25888 39313 25891
rect 38712 25860 39313 25888
rect 38712 25848 38718 25860
rect 39301 25857 39313 25860
rect 39347 25857 39359 25891
rect 39301 25851 39359 25857
rect 39669 25891 39727 25897
rect 39669 25857 39681 25891
rect 39715 25888 39727 25891
rect 40218 25888 40224 25900
rect 39715 25860 40224 25888
rect 39715 25857 39727 25860
rect 39669 25851 39727 25857
rect 40218 25848 40224 25860
rect 40276 25848 40282 25900
rect 40494 25848 40500 25900
rect 40552 25888 40558 25900
rect 41049 25891 41107 25897
rect 41049 25888 41061 25891
rect 40552 25860 41061 25888
rect 40552 25848 40558 25860
rect 41049 25857 41061 25860
rect 41095 25857 41107 25891
rect 41049 25851 41107 25857
rect 41138 25848 41144 25900
rect 41196 25888 41202 25900
rect 41966 25888 41972 25900
rect 41196 25860 41972 25888
rect 41196 25848 41202 25860
rect 41966 25848 41972 25860
rect 42024 25848 42030 25900
rect 42613 25891 42671 25897
rect 42613 25857 42625 25891
rect 42659 25888 42671 25891
rect 42978 25888 42984 25900
rect 42659 25860 42984 25888
rect 42659 25857 42671 25860
rect 42613 25851 42671 25857
rect 42978 25848 42984 25860
rect 43036 25848 43042 25900
rect 43717 25891 43775 25897
rect 43717 25857 43729 25891
rect 43763 25888 43775 25891
rect 43990 25888 43996 25900
rect 43763 25860 43996 25888
rect 43763 25857 43775 25860
rect 43717 25851 43775 25857
rect 43990 25848 43996 25860
rect 44048 25848 44054 25900
rect 44453 25891 44511 25897
rect 44453 25857 44465 25891
rect 44499 25888 44511 25891
rect 45830 25888 45836 25900
rect 44499 25860 45836 25888
rect 44499 25857 44511 25860
rect 44453 25851 44511 25857
rect 45830 25848 45836 25860
rect 45888 25848 45894 25900
rect 46014 25848 46020 25900
rect 46072 25888 46078 25900
rect 46124 25897 46152 25928
rect 47118 25916 47124 25928
rect 47176 25916 47182 25968
rect 47578 25916 47584 25968
rect 47636 25956 47642 25968
rect 49068 25965 49096 25996
rect 49510 25984 49516 25996
rect 49568 26024 49574 26036
rect 49697 26027 49755 26033
rect 49697 26024 49709 26027
rect 49568 25996 49709 26024
rect 49568 25984 49574 25996
rect 49697 25993 49709 25996
rect 49743 25993 49755 26027
rect 49697 25987 49755 25993
rect 50433 26027 50491 26033
rect 50433 25993 50445 26027
rect 50479 26024 50491 26027
rect 50982 26024 50988 26036
rect 50479 25996 50988 26024
rect 50479 25993 50491 25996
rect 50433 25987 50491 25993
rect 50982 25984 50988 25996
rect 51040 25984 51046 26036
rect 52089 26027 52147 26033
rect 52089 25993 52101 26027
rect 52135 26024 52147 26027
rect 52362 26024 52368 26036
rect 52135 25996 52368 26024
rect 52135 25993 52147 25996
rect 52089 25987 52147 25993
rect 52362 25984 52368 25996
rect 52420 25984 52426 26036
rect 53653 26027 53711 26033
rect 53653 25993 53665 26027
rect 53699 26024 53711 26027
rect 54570 26024 54576 26036
rect 53699 25996 54576 26024
rect 53699 25993 53711 25996
rect 53653 25987 53711 25993
rect 54570 25984 54576 25996
rect 54628 26024 54634 26036
rect 55677 26027 55735 26033
rect 55677 26024 55689 26027
rect 54628 25996 55689 26024
rect 54628 25984 54634 25996
rect 55677 25993 55689 25996
rect 55723 25993 55735 26027
rect 55677 25987 55735 25993
rect 56134 25984 56140 26036
rect 56192 26024 56198 26036
rect 56229 26027 56287 26033
rect 56229 26024 56241 26027
rect 56192 25996 56241 26024
rect 56192 25984 56198 25996
rect 56229 25993 56241 25996
rect 56275 26024 56287 26027
rect 58250 26024 58256 26036
rect 56275 25996 58256 26024
rect 56275 25993 56287 25996
rect 56229 25987 56287 25993
rect 58250 25984 58256 25996
rect 58308 25984 58314 26036
rect 48041 25959 48099 25965
rect 48041 25956 48053 25959
rect 47636 25928 48053 25956
rect 47636 25916 47642 25928
rect 48041 25925 48053 25928
rect 48087 25925 48099 25959
rect 48041 25919 48099 25925
rect 49053 25959 49111 25965
rect 49053 25925 49065 25959
rect 49099 25925 49111 25959
rect 49053 25919 49111 25925
rect 49237 25959 49295 25965
rect 49237 25925 49249 25959
rect 49283 25956 49295 25959
rect 50154 25956 50160 25968
rect 49283 25928 50160 25956
rect 49283 25925 49295 25928
rect 49237 25919 49295 25925
rect 46109 25891 46167 25897
rect 46109 25888 46121 25891
rect 46072 25860 46121 25888
rect 46072 25848 46078 25860
rect 46109 25857 46121 25860
rect 46155 25857 46167 25891
rect 46109 25851 46167 25857
rect 47026 25848 47032 25900
rect 47084 25888 47090 25900
rect 47949 25891 48007 25897
rect 47949 25888 47961 25891
rect 47084 25860 47961 25888
rect 47084 25848 47090 25860
rect 47949 25857 47961 25860
rect 47995 25857 48007 25891
rect 47949 25851 48007 25857
rect 48133 25891 48191 25897
rect 48133 25857 48145 25891
rect 48179 25888 48191 25891
rect 48222 25888 48228 25900
rect 48179 25860 48228 25888
rect 48179 25857 48191 25860
rect 48133 25851 48191 25857
rect 48222 25848 48228 25860
rect 48280 25848 48286 25900
rect 48317 25891 48375 25897
rect 48317 25857 48329 25891
rect 48363 25857 48375 25891
rect 48317 25851 48375 25857
rect 39209 25823 39267 25829
rect 39209 25789 39221 25823
rect 39255 25820 39267 25823
rect 39850 25820 39856 25832
rect 39255 25792 39856 25820
rect 39255 25789 39267 25792
rect 39209 25783 39267 25789
rect 39850 25780 39856 25792
rect 39908 25780 39914 25832
rect 45922 25820 45928 25832
rect 45883 25792 45928 25820
rect 45922 25780 45928 25792
rect 45980 25780 45986 25832
rect 48332 25820 48360 25851
rect 48406 25848 48412 25900
rect 48464 25888 48470 25900
rect 49252 25888 49280 25919
rect 50154 25916 50160 25928
rect 50212 25916 50218 25968
rect 50798 25916 50804 25968
rect 50856 25956 50862 25968
rect 50893 25959 50951 25965
rect 50893 25956 50905 25959
rect 50856 25928 50905 25956
rect 50856 25916 50862 25928
rect 50893 25925 50905 25928
rect 50939 25925 50951 25959
rect 50893 25919 50951 25925
rect 55217 25959 55275 25965
rect 55217 25925 55229 25959
rect 55263 25956 55275 25959
rect 56152 25956 56180 25984
rect 55263 25928 56180 25956
rect 55263 25925 55275 25928
rect 55217 25919 55275 25925
rect 48464 25860 49280 25888
rect 49697 25891 49755 25897
rect 48464 25848 48470 25860
rect 49697 25857 49709 25891
rect 49743 25888 49755 25891
rect 49786 25888 49792 25900
rect 49743 25860 49792 25888
rect 49743 25857 49755 25860
rect 49697 25851 49755 25857
rect 49786 25848 49792 25860
rect 49844 25848 49850 25900
rect 49878 25848 49884 25900
rect 49936 25888 49942 25900
rect 49936 25860 49981 25888
rect 49936 25848 49942 25860
rect 48332 25792 51580 25820
rect 40034 25752 40040 25764
rect 38580 25724 40040 25752
rect 40034 25712 40040 25724
rect 40092 25712 40098 25764
rect 47854 25712 47860 25764
rect 47912 25752 47918 25764
rect 50798 25752 50804 25764
rect 47912 25724 50804 25752
rect 47912 25712 47918 25724
rect 50798 25712 50804 25724
rect 50856 25712 50862 25764
rect 51552 25696 51580 25792
rect 38473 25687 38531 25693
rect 38473 25653 38485 25687
rect 38519 25684 38531 25687
rect 38930 25684 38936 25696
rect 38519 25656 38936 25684
rect 38519 25653 38531 25656
rect 38473 25647 38531 25653
rect 38930 25644 38936 25656
rect 38988 25644 38994 25696
rect 44174 25644 44180 25696
rect 44232 25684 44238 25696
rect 44269 25687 44327 25693
rect 44269 25684 44281 25687
rect 44232 25656 44281 25684
rect 44232 25644 44238 25656
rect 44269 25653 44281 25656
rect 44315 25653 44327 25687
rect 44269 25647 44327 25653
rect 44358 25644 44364 25696
rect 44416 25684 44422 25696
rect 44910 25684 44916 25696
rect 44416 25656 44916 25684
rect 44416 25644 44422 25656
rect 44910 25644 44916 25656
rect 44968 25644 44974 25696
rect 47765 25687 47823 25693
rect 47765 25653 47777 25687
rect 47811 25684 47823 25687
rect 48682 25684 48688 25696
rect 47811 25656 48688 25684
rect 47811 25653 47823 25656
rect 47765 25647 47823 25653
rect 48682 25644 48688 25656
rect 48740 25644 48746 25696
rect 48866 25684 48872 25696
rect 48827 25656 48872 25684
rect 48866 25644 48872 25656
rect 48924 25644 48930 25696
rect 51534 25684 51540 25696
rect 51495 25656 51540 25684
rect 51534 25644 51540 25656
rect 51592 25644 51598 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 35529 25483 35587 25489
rect 35529 25449 35541 25483
rect 35575 25480 35587 25483
rect 36170 25480 36176 25492
rect 35575 25452 36176 25480
rect 35575 25449 35587 25452
rect 35529 25443 35587 25449
rect 36170 25440 36176 25452
rect 36228 25440 36234 25492
rect 37458 25480 37464 25492
rect 37419 25452 37464 25480
rect 37458 25440 37464 25452
rect 37516 25440 37522 25492
rect 38010 25480 38016 25492
rect 37971 25452 38016 25480
rect 38010 25440 38016 25452
rect 38068 25440 38074 25492
rect 38102 25440 38108 25492
rect 38160 25480 38166 25492
rect 39114 25480 39120 25492
rect 38160 25452 39120 25480
rect 38160 25440 38166 25452
rect 39114 25440 39120 25452
rect 39172 25440 39178 25492
rect 39301 25483 39359 25489
rect 39301 25449 39313 25483
rect 39347 25480 39359 25483
rect 40126 25480 40132 25492
rect 39347 25452 40132 25480
rect 39347 25449 39359 25452
rect 39301 25443 39359 25449
rect 40126 25440 40132 25452
rect 40184 25440 40190 25492
rect 40494 25480 40500 25492
rect 40455 25452 40500 25480
rect 40494 25440 40500 25452
rect 40552 25440 40558 25492
rect 41138 25440 41144 25492
rect 41196 25440 41202 25492
rect 43070 25440 43076 25492
rect 43128 25480 43134 25492
rect 43441 25483 43499 25489
rect 43441 25480 43453 25483
rect 43128 25452 43453 25480
rect 43128 25440 43134 25452
rect 43441 25449 43453 25452
rect 43487 25449 43499 25483
rect 43441 25443 43499 25449
rect 43806 25440 43812 25492
rect 43864 25480 43870 25492
rect 43993 25483 44051 25489
rect 43993 25480 44005 25483
rect 43864 25452 44005 25480
rect 43864 25440 43870 25452
rect 43993 25449 44005 25452
rect 44039 25480 44051 25483
rect 44545 25483 44603 25489
rect 44545 25480 44557 25483
rect 44039 25452 44557 25480
rect 44039 25449 44051 25452
rect 43993 25443 44051 25449
rect 44545 25449 44557 25452
rect 44591 25449 44603 25483
rect 44545 25443 44603 25449
rect 46290 25440 46296 25492
rect 46348 25480 46354 25492
rect 47302 25480 47308 25492
rect 46348 25452 47308 25480
rect 46348 25440 46354 25452
rect 47302 25440 47308 25452
rect 47360 25440 47366 25492
rect 48222 25480 48228 25492
rect 48183 25452 48228 25480
rect 48222 25440 48228 25452
rect 48280 25440 48286 25492
rect 49050 25480 49056 25492
rect 49011 25452 49056 25480
rect 49050 25440 49056 25452
rect 49108 25440 49114 25492
rect 52178 25480 52184 25492
rect 51046 25452 52184 25480
rect 37642 25304 37648 25356
rect 37700 25344 37706 25356
rect 38028 25344 38056 25440
rect 38381 25415 38439 25421
rect 38381 25381 38393 25415
rect 38427 25412 38439 25415
rect 39850 25412 39856 25424
rect 38427 25384 39856 25412
rect 38427 25381 38439 25384
rect 38381 25375 38439 25381
rect 39850 25372 39856 25384
rect 39908 25372 39914 25424
rect 41156 25412 41184 25440
rect 40972 25384 41184 25412
rect 42889 25415 42947 25421
rect 40402 25344 40408 25356
rect 37700 25316 37780 25344
rect 38028 25316 38976 25344
rect 37700 25304 37706 25316
rect 31754 25236 31760 25288
rect 31812 25276 31818 25288
rect 34333 25279 34391 25285
rect 34333 25276 34345 25279
rect 31812 25248 34345 25276
rect 31812 25236 31818 25248
rect 34333 25245 34345 25248
rect 34379 25276 34391 25279
rect 35437 25279 35495 25285
rect 35437 25276 35449 25279
rect 34379 25248 35449 25276
rect 34379 25245 34391 25248
rect 34333 25239 34391 25245
rect 35437 25245 35449 25248
rect 35483 25245 35495 25279
rect 36446 25276 36452 25288
rect 36407 25248 36452 25276
rect 35437 25239 35495 25245
rect 34790 25100 34796 25152
rect 34848 25140 34854 25152
rect 34885 25143 34943 25149
rect 34885 25140 34897 25143
rect 34848 25112 34897 25140
rect 34848 25100 34854 25112
rect 34885 25109 34897 25112
rect 34931 25109 34943 25143
rect 35452 25140 35480 25239
rect 36446 25236 36452 25248
rect 36504 25236 36510 25288
rect 36998 25236 37004 25288
rect 37056 25276 37062 25288
rect 37752 25276 37780 25316
rect 38194 25276 38200 25288
rect 37056 25248 37688 25276
rect 37752 25248 38200 25276
rect 37056 25236 37062 25248
rect 36265 25211 36323 25217
rect 36265 25177 36277 25211
rect 36311 25208 36323 25211
rect 36538 25208 36544 25220
rect 36311 25180 36544 25208
rect 36311 25177 36323 25180
rect 36265 25171 36323 25177
rect 36538 25168 36544 25180
rect 36596 25168 36602 25220
rect 36633 25211 36691 25217
rect 36633 25177 36645 25211
rect 36679 25208 36691 25211
rect 37185 25211 37243 25217
rect 37185 25208 37197 25211
rect 36679 25180 37197 25208
rect 36679 25177 36691 25180
rect 36633 25171 36691 25177
rect 37185 25177 37197 25180
rect 37231 25177 37243 25211
rect 37660 25208 37688 25248
rect 38194 25236 38200 25248
rect 38252 25236 38258 25288
rect 38470 25276 38476 25288
rect 38431 25248 38476 25276
rect 38470 25236 38476 25248
rect 38528 25236 38534 25288
rect 38948 25285 38976 25316
rect 39224 25316 40408 25344
rect 38933 25279 38991 25285
rect 38933 25245 38945 25279
rect 38979 25245 38991 25279
rect 38933 25239 38991 25245
rect 39022 25236 39028 25288
rect 39080 25276 39086 25288
rect 39080 25248 39125 25276
rect 39080 25236 39086 25248
rect 38838 25208 38844 25220
rect 37660 25180 38844 25208
rect 37185 25171 37243 25177
rect 38838 25168 38844 25180
rect 38896 25208 38902 25220
rect 39224 25208 39252 25316
rect 40402 25304 40408 25316
rect 40460 25304 40466 25356
rect 40589 25347 40647 25353
rect 40589 25313 40601 25347
rect 40635 25344 40647 25347
rect 40862 25344 40868 25356
rect 40635 25316 40868 25344
rect 40635 25313 40647 25316
rect 40589 25307 40647 25313
rect 40862 25304 40868 25316
rect 40920 25304 40926 25356
rect 40681 25279 40739 25285
rect 40681 25245 40693 25279
rect 40727 25276 40739 25279
rect 40972 25276 41000 25384
rect 42889 25381 42901 25415
rect 42935 25412 42947 25415
rect 43162 25412 43168 25424
rect 42935 25384 43168 25412
rect 42935 25381 42947 25384
rect 42889 25375 42947 25381
rect 43162 25372 43168 25384
rect 43220 25372 43226 25424
rect 46474 25412 46480 25424
rect 46387 25384 46480 25412
rect 46474 25372 46480 25384
rect 46532 25412 46538 25424
rect 47489 25415 47547 25421
rect 47489 25412 47501 25415
rect 46532 25384 47501 25412
rect 46532 25372 46538 25384
rect 47489 25381 47501 25384
rect 47535 25412 47547 25415
rect 48406 25412 48412 25424
rect 47535 25384 48412 25412
rect 47535 25381 47547 25384
rect 47489 25375 47547 25381
rect 48406 25372 48412 25384
rect 48464 25372 48470 25424
rect 51046 25412 51074 25452
rect 52178 25440 52184 25452
rect 52236 25480 52242 25492
rect 54389 25483 54447 25489
rect 54389 25480 54401 25483
rect 52236 25452 54401 25480
rect 52236 25440 52242 25452
rect 54389 25449 54401 25452
rect 54435 25449 54447 25483
rect 54389 25443 54447 25449
rect 52638 25412 52644 25424
rect 49896 25384 51074 25412
rect 52551 25384 52644 25412
rect 41141 25347 41199 25353
rect 41141 25313 41153 25347
rect 41187 25344 41199 25347
rect 42702 25344 42708 25356
rect 41187 25316 42708 25344
rect 41187 25313 41199 25316
rect 41141 25307 41199 25313
rect 42702 25304 42708 25316
rect 42760 25304 42766 25356
rect 40727 25248 41000 25276
rect 40727 25245 40739 25248
rect 40681 25239 40739 25245
rect 45094 25236 45100 25288
rect 45152 25276 45158 25288
rect 45189 25279 45247 25285
rect 45189 25276 45201 25279
rect 45152 25248 45201 25276
rect 45152 25236 45158 25248
rect 45189 25245 45201 25248
rect 45235 25245 45247 25279
rect 45189 25239 45247 25245
rect 46198 25236 46204 25288
rect 46256 25276 46262 25288
rect 46492 25285 46520 25372
rect 49896 25356 49924 25384
rect 52638 25372 52644 25384
rect 52696 25412 52702 25424
rect 57974 25412 57980 25424
rect 52696 25384 57980 25412
rect 52696 25372 52702 25384
rect 57974 25372 57980 25384
rect 58032 25372 58038 25424
rect 47121 25347 47179 25353
rect 47121 25313 47133 25347
rect 47167 25344 47179 25347
rect 49697 25347 49755 25353
rect 47167 25316 48360 25344
rect 47167 25313 47179 25316
rect 47121 25307 47179 25313
rect 48332 25288 48360 25316
rect 49697 25313 49709 25347
rect 49743 25344 49755 25347
rect 49878 25344 49884 25356
rect 49743 25316 49884 25344
rect 49743 25313 49755 25316
rect 49697 25307 49755 25313
rect 49878 25304 49884 25316
rect 49936 25304 49942 25356
rect 50062 25304 50068 25356
rect 50120 25344 50126 25356
rect 50120 25316 50844 25344
rect 50120 25304 50126 25316
rect 46293 25279 46351 25285
rect 46293 25276 46305 25279
rect 46256 25248 46305 25276
rect 46256 25236 46262 25248
rect 46293 25245 46305 25248
rect 46339 25245 46351 25279
rect 46293 25239 46351 25245
rect 46477 25279 46535 25285
rect 46477 25245 46489 25279
rect 46523 25245 46535 25279
rect 47026 25276 47032 25288
rect 46987 25248 47032 25276
rect 46477 25239 46535 25245
rect 47026 25236 47032 25248
rect 47084 25236 47090 25288
rect 47210 25276 47216 25288
rect 47171 25248 47216 25276
rect 47210 25236 47216 25248
rect 47268 25236 47274 25288
rect 47302 25236 47308 25288
rect 47360 25276 47366 25288
rect 48314 25276 48320 25288
rect 47360 25248 47405 25276
rect 48275 25248 48320 25276
rect 47360 25236 47366 25248
rect 48314 25236 48320 25248
rect 48372 25236 48378 25288
rect 48869 25279 48927 25285
rect 48869 25245 48881 25279
rect 48915 25245 48927 25279
rect 48869 25239 48927 25245
rect 49145 25279 49203 25285
rect 49145 25245 49157 25279
rect 49191 25276 49203 25279
rect 49602 25276 49608 25288
rect 49191 25248 49608 25276
rect 49191 25245 49203 25248
rect 49145 25239 49203 25245
rect 38896 25180 39252 25208
rect 39408 25180 40448 25208
rect 38896 25168 38902 25180
rect 39408 25140 39436 25180
rect 35452 25112 39436 25140
rect 34885 25103 34943 25109
rect 39850 25100 39856 25152
rect 39908 25140 39914 25152
rect 40310 25140 40316 25152
rect 39908 25112 40316 25140
rect 39908 25100 39914 25112
rect 40310 25100 40316 25112
rect 40368 25100 40374 25152
rect 40420 25140 40448 25180
rect 41046 25168 41052 25220
rect 41104 25208 41110 25220
rect 41417 25211 41475 25217
rect 41417 25208 41429 25211
rect 41104 25180 41429 25208
rect 41104 25168 41110 25180
rect 41417 25177 41429 25180
rect 41463 25177 41475 25211
rect 43070 25208 43076 25220
rect 42642 25180 43076 25208
rect 41417 25171 41475 25177
rect 43070 25168 43076 25180
rect 43128 25168 43134 25220
rect 46934 25168 46940 25220
rect 46992 25208 46998 25220
rect 48884 25208 48912 25239
rect 49602 25236 49608 25248
rect 49660 25236 49666 25288
rect 50154 25236 50160 25288
rect 50212 25276 50218 25288
rect 50816 25285 50844 25316
rect 51074 25304 51080 25356
rect 51132 25344 51138 25356
rect 51261 25347 51319 25353
rect 51261 25344 51273 25347
rect 51132 25316 51273 25344
rect 51132 25304 51138 25316
rect 51261 25313 51273 25316
rect 51307 25313 51319 25347
rect 51261 25307 51319 25313
rect 50617 25279 50675 25285
rect 50617 25276 50629 25279
rect 50212 25248 50629 25276
rect 50212 25236 50218 25248
rect 50617 25245 50629 25248
rect 50663 25245 50675 25279
rect 50617 25239 50675 25245
rect 50801 25279 50859 25285
rect 50801 25245 50813 25279
rect 50847 25276 50859 25279
rect 50982 25276 50988 25288
rect 50847 25248 50988 25276
rect 50847 25245 50859 25248
rect 50801 25239 50859 25245
rect 50982 25236 50988 25248
rect 51040 25236 51046 25288
rect 51276 25276 51304 25307
rect 51810 25276 51816 25288
rect 51276 25248 51816 25276
rect 51810 25236 51816 25248
rect 51868 25236 51874 25288
rect 46992 25180 48912 25208
rect 48961 25211 49019 25217
rect 46992 25168 46998 25180
rect 48961 25177 48973 25211
rect 49007 25208 49019 25211
rect 49694 25208 49700 25220
rect 49007 25180 49700 25208
rect 49007 25177 49019 25180
rect 48961 25171 49019 25177
rect 42242 25140 42248 25152
rect 40420 25112 42248 25140
rect 42242 25100 42248 25112
rect 42300 25100 42306 25152
rect 45186 25100 45192 25152
rect 45244 25140 45250 25152
rect 45281 25143 45339 25149
rect 45281 25140 45293 25143
rect 45244 25112 45293 25140
rect 45244 25100 45250 25112
rect 45281 25109 45293 25112
rect 45327 25109 45339 25143
rect 46290 25140 46296 25152
rect 46251 25112 46296 25140
rect 45281 25103 45339 25109
rect 46290 25100 46296 25112
rect 46348 25100 46354 25152
rect 47578 25100 47584 25152
rect 47636 25140 47642 25152
rect 48222 25140 48228 25152
rect 47636 25112 48228 25140
rect 47636 25100 47642 25112
rect 48222 25100 48228 25112
rect 48280 25140 48286 25152
rect 48976 25140 49004 25171
rect 49694 25168 49700 25180
rect 49752 25168 49758 25220
rect 51074 25168 51080 25220
rect 51132 25208 51138 25220
rect 51506 25211 51564 25217
rect 51506 25208 51518 25211
rect 51132 25180 51518 25208
rect 51132 25168 51138 25180
rect 51506 25177 51518 25180
rect 51552 25177 51564 25211
rect 51506 25171 51564 25177
rect 48280 25112 49004 25140
rect 50709 25143 50767 25149
rect 48280 25100 48286 25112
rect 50709 25109 50721 25143
rect 50755 25140 50767 25143
rect 51626 25140 51632 25152
rect 50755 25112 51632 25140
rect 50755 25109 50767 25112
rect 50709 25103 50767 25109
rect 51626 25100 51632 25112
rect 51684 25100 51690 25152
rect 1104 25050 58880 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 58880 25050
rect 1104 24976 58880 24998
rect 36357 24939 36415 24945
rect 36357 24905 36369 24939
rect 36403 24936 36415 24939
rect 36446 24936 36452 24948
rect 36403 24908 36452 24936
rect 36403 24905 36415 24908
rect 36357 24899 36415 24905
rect 36446 24896 36452 24908
rect 36504 24896 36510 24948
rect 37550 24896 37556 24948
rect 37608 24936 37614 24948
rect 40126 24936 40132 24948
rect 37608 24908 37780 24936
rect 37608 24896 37614 24908
rect 34606 24800 34612 24812
rect 34567 24772 34612 24800
rect 34606 24760 34612 24772
rect 34664 24760 34670 24812
rect 35986 24760 35992 24812
rect 36044 24760 36050 24812
rect 36464 24800 36492 24896
rect 37458 24828 37464 24880
rect 37516 24868 37522 24880
rect 37752 24877 37780 24908
rect 39316 24908 40132 24936
rect 37737 24871 37795 24877
rect 37516 24840 37688 24868
rect 37516 24828 37522 24840
rect 37660 24809 37688 24840
rect 37737 24837 37749 24871
rect 37783 24837 37795 24871
rect 38838 24868 38844 24880
rect 38799 24840 38844 24868
rect 37737 24831 37795 24837
rect 38838 24828 38844 24840
rect 38896 24828 38902 24880
rect 37645 24803 37703 24809
rect 36464 24772 37596 24800
rect 34885 24735 34943 24741
rect 34885 24701 34897 24735
rect 34931 24732 34943 24735
rect 37461 24735 37519 24741
rect 37461 24732 37473 24735
rect 34931 24704 37473 24732
rect 34931 24701 34943 24704
rect 34885 24695 34943 24701
rect 37461 24701 37473 24704
rect 37507 24701 37519 24735
rect 37568 24732 37596 24772
rect 37645 24769 37657 24803
rect 37691 24769 37703 24803
rect 37645 24763 37703 24769
rect 37826 24760 37832 24812
rect 37884 24800 37890 24812
rect 37967 24803 38025 24809
rect 37884 24772 37929 24800
rect 37884 24760 37890 24772
rect 37967 24769 37979 24803
rect 38013 24800 38025 24803
rect 38930 24800 38936 24812
rect 38013 24772 38332 24800
rect 38891 24772 38936 24800
rect 38013 24769 38025 24772
rect 37967 24763 38025 24769
rect 38105 24735 38163 24741
rect 38105 24732 38117 24735
rect 37568 24704 38117 24732
rect 37461 24695 37519 24701
rect 38105 24701 38117 24704
rect 38151 24701 38163 24735
rect 38304 24732 38332 24772
rect 38930 24760 38936 24772
rect 38988 24760 38994 24812
rect 39209 24803 39267 24809
rect 39209 24769 39221 24803
rect 39255 24800 39267 24803
rect 39316 24800 39344 24908
rect 40126 24896 40132 24908
rect 40184 24896 40190 24948
rect 40862 24896 40868 24948
rect 40920 24936 40926 24948
rect 40920 24908 41920 24936
rect 40920 24896 40926 24908
rect 39837 24871 39895 24877
rect 39837 24837 39849 24871
rect 39883 24868 39895 24871
rect 40034 24868 40040 24880
rect 39883 24837 39896 24868
rect 39995 24840 40040 24868
rect 39837 24831 39896 24837
rect 39255 24772 39344 24800
rect 39255 24769 39267 24772
rect 39209 24763 39267 24769
rect 39390 24760 39396 24812
rect 39448 24800 39454 24812
rect 39868 24800 39896 24831
rect 40034 24828 40040 24840
rect 40092 24828 40098 24880
rect 40310 24828 40316 24880
rect 40368 24868 40374 24880
rect 41598 24868 41604 24880
rect 40368 24840 41604 24868
rect 40368 24828 40374 24840
rect 41598 24828 41604 24840
rect 41656 24828 41662 24880
rect 41785 24871 41843 24877
rect 41785 24837 41797 24871
rect 41831 24837 41843 24871
rect 41785 24831 41843 24837
rect 39448 24772 39896 24800
rect 39448 24760 39454 24772
rect 38838 24732 38844 24744
rect 38304 24704 38844 24732
rect 38105 24695 38163 24701
rect 38120 24664 38148 24695
rect 38838 24692 38844 24704
rect 38896 24692 38902 24744
rect 38286 24664 38292 24676
rect 38120 24636 38292 24664
rect 38286 24624 38292 24636
rect 38344 24624 38350 24676
rect 39666 24664 39672 24676
rect 39627 24636 39672 24664
rect 39666 24624 39672 24636
rect 39724 24624 39730 24676
rect 39868 24664 39896 24772
rect 40402 24760 40408 24812
rect 40460 24800 40466 24812
rect 40681 24803 40739 24809
rect 40681 24800 40693 24803
rect 40460 24772 40693 24800
rect 40460 24760 40466 24772
rect 40681 24769 40693 24772
rect 40727 24769 40739 24803
rect 40862 24800 40868 24812
rect 40823 24772 40868 24800
rect 40681 24763 40739 24769
rect 40862 24760 40868 24772
rect 40920 24760 40926 24812
rect 40954 24760 40960 24812
rect 41012 24800 41018 24812
rect 41509 24803 41567 24809
rect 41509 24800 41521 24803
rect 41012 24772 41521 24800
rect 41012 24760 41018 24772
rect 41509 24769 41521 24772
rect 41555 24769 41567 24803
rect 41800 24800 41828 24831
rect 41509 24763 41567 24769
rect 41616 24772 41828 24800
rect 39942 24692 39948 24744
rect 40000 24732 40006 24744
rect 41616 24732 41644 24772
rect 41782 24732 41788 24744
rect 40000 24704 41644 24732
rect 41743 24704 41788 24732
rect 40000 24692 40006 24704
rect 41782 24692 41788 24704
rect 41840 24692 41846 24744
rect 41892 24732 41920 24908
rect 45833 24871 45891 24877
rect 45833 24837 45845 24871
rect 45879 24868 45891 24871
rect 45922 24868 45928 24880
rect 45879 24840 45928 24868
rect 45879 24837 45891 24840
rect 45833 24831 45891 24837
rect 45922 24828 45928 24840
rect 45980 24828 45986 24880
rect 41966 24760 41972 24812
rect 42024 24800 42030 24812
rect 42797 24803 42855 24809
rect 42797 24800 42809 24803
rect 42024 24772 42809 24800
rect 42024 24760 42030 24772
rect 42797 24769 42809 24772
rect 42843 24769 42855 24803
rect 42797 24763 42855 24769
rect 42886 24760 42892 24812
rect 42944 24800 42950 24812
rect 42944 24772 42989 24800
rect 42944 24760 42950 24772
rect 45186 24760 45192 24812
rect 45244 24760 45250 24812
rect 45370 24760 45376 24812
rect 45428 24800 45434 24812
rect 46477 24803 46535 24809
rect 46477 24800 46489 24803
rect 45428 24772 46489 24800
rect 45428 24760 45434 24772
rect 46477 24769 46489 24772
rect 46523 24769 46535 24803
rect 46477 24763 46535 24769
rect 46661 24803 46719 24809
rect 46661 24769 46673 24803
rect 46707 24800 46719 24803
rect 46934 24800 46940 24812
rect 46707 24772 46940 24800
rect 46707 24769 46719 24772
rect 46661 24763 46719 24769
rect 46934 24760 46940 24772
rect 46992 24760 46998 24812
rect 47854 24800 47860 24812
rect 47815 24772 47860 24800
rect 47854 24760 47860 24772
rect 47912 24760 47918 24812
rect 48774 24800 48780 24812
rect 48735 24772 48780 24800
rect 48774 24760 48780 24772
rect 48832 24760 48838 24812
rect 51166 24800 51172 24812
rect 51127 24772 51172 24800
rect 51166 24760 51172 24772
rect 51224 24760 51230 24812
rect 51261 24803 51319 24809
rect 51261 24769 51273 24803
rect 51307 24769 51319 24803
rect 51261 24763 51319 24769
rect 51537 24803 51595 24809
rect 51537 24769 51549 24803
rect 51583 24800 51595 24803
rect 52638 24800 52644 24812
rect 51583 24772 52644 24800
rect 51583 24769 51595 24772
rect 51537 24763 51595 24769
rect 42613 24735 42671 24741
rect 42613 24732 42625 24735
rect 41892 24704 42625 24732
rect 42613 24701 42625 24704
rect 42659 24701 42671 24735
rect 42613 24695 42671 24701
rect 42702 24692 42708 24744
rect 42760 24732 42766 24744
rect 43809 24735 43867 24741
rect 43809 24732 43821 24735
rect 42760 24704 43821 24732
rect 42760 24692 42766 24704
rect 43809 24701 43821 24704
rect 43855 24701 43867 24735
rect 43809 24695 43867 24701
rect 44085 24735 44143 24741
rect 44085 24701 44097 24735
rect 44131 24732 44143 24735
rect 44174 24732 44180 24744
rect 44131 24704 44180 24732
rect 44131 24701 44143 24704
rect 44085 24695 44143 24701
rect 44174 24692 44180 24704
rect 44232 24692 44238 24744
rect 50985 24735 51043 24741
rect 50985 24701 50997 24735
rect 51031 24732 51043 24735
rect 51074 24732 51080 24744
rect 51031 24704 51080 24732
rect 51031 24701 51043 24704
rect 50985 24695 51043 24701
rect 51074 24692 51080 24704
rect 51132 24692 51138 24744
rect 39868 24636 40264 24664
rect 37550 24556 37556 24608
rect 37608 24596 37614 24608
rect 39022 24596 39028 24608
rect 37608 24568 39028 24596
rect 37608 24556 37614 24568
rect 39022 24556 39028 24568
rect 39080 24556 39086 24608
rect 39298 24556 39304 24608
rect 39356 24596 39362 24608
rect 39850 24596 39856 24608
rect 39356 24568 39856 24596
rect 39356 24556 39362 24568
rect 39850 24556 39856 24568
rect 39908 24556 39914 24608
rect 40236 24596 40264 24636
rect 41046 24624 41052 24676
rect 41104 24664 41110 24676
rect 46845 24667 46903 24673
rect 41104 24636 41149 24664
rect 41524 24636 42748 24664
rect 41104 24624 41110 24636
rect 41524 24596 41552 24636
rect 40236 24568 41552 24596
rect 41598 24556 41604 24608
rect 41656 24596 41662 24608
rect 42720 24605 42748 24636
rect 46845 24633 46857 24667
rect 46891 24664 46903 24667
rect 47026 24664 47032 24676
rect 46891 24636 47032 24664
rect 46891 24633 46903 24636
rect 46845 24627 46903 24633
rect 47026 24624 47032 24636
rect 47084 24624 47090 24676
rect 48682 24624 48688 24676
rect 48740 24664 48746 24676
rect 51276 24664 51304 24763
rect 52638 24760 52644 24772
rect 52696 24760 52702 24812
rect 51445 24735 51503 24741
rect 51445 24701 51457 24735
rect 51491 24732 51503 24735
rect 51626 24732 51632 24744
rect 51491 24704 51632 24732
rect 51491 24701 51503 24704
rect 51445 24695 51503 24701
rect 51626 24692 51632 24704
rect 51684 24692 51690 24744
rect 48740 24636 51304 24664
rect 48740 24624 48746 24636
rect 42705 24599 42763 24605
rect 41656 24568 41701 24596
rect 41656 24556 41662 24568
rect 42705 24565 42717 24599
rect 42751 24565 42763 24599
rect 42705 24559 42763 24565
rect 46661 24599 46719 24605
rect 46661 24565 46673 24599
rect 46707 24596 46719 24599
rect 47578 24596 47584 24608
rect 46707 24568 47584 24596
rect 46707 24565 46719 24568
rect 46661 24559 46719 24565
rect 47578 24556 47584 24568
rect 47636 24556 47642 24608
rect 50246 24596 50252 24608
rect 50207 24568 50252 24596
rect 50246 24556 50252 24568
rect 50304 24556 50310 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 35805 24395 35863 24401
rect 35805 24361 35817 24395
rect 35851 24392 35863 24395
rect 35986 24392 35992 24404
rect 35851 24364 35992 24392
rect 35851 24361 35863 24364
rect 35805 24355 35863 24361
rect 35986 24352 35992 24364
rect 36044 24352 36050 24404
rect 40770 24352 40776 24404
rect 40828 24392 40834 24404
rect 42797 24395 42855 24401
rect 42797 24392 42809 24395
rect 40828 24364 42809 24392
rect 40828 24352 40834 24364
rect 42797 24361 42809 24364
rect 42843 24361 42855 24395
rect 42797 24355 42855 24361
rect 43070 24352 43076 24404
rect 43128 24392 43134 24404
rect 43441 24395 43499 24401
rect 43441 24392 43453 24395
rect 43128 24364 43453 24392
rect 43128 24352 43134 24364
rect 43441 24361 43453 24364
rect 43487 24361 43499 24395
rect 43441 24355 43499 24361
rect 44085 24395 44143 24401
rect 44085 24361 44097 24395
rect 44131 24392 44143 24395
rect 44910 24392 44916 24404
rect 44131 24364 44916 24392
rect 44131 24361 44143 24364
rect 44085 24355 44143 24361
rect 44910 24352 44916 24364
rect 44968 24352 44974 24404
rect 46477 24395 46535 24401
rect 46477 24361 46489 24395
rect 46523 24392 46535 24395
rect 47026 24392 47032 24404
rect 46523 24364 47032 24392
rect 46523 24361 46535 24364
rect 46477 24355 46535 24361
rect 47026 24352 47032 24364
rect 47084 24352 47090 24404
rect 48314 24352 48320 24404
rect 48372 24392 48378 24404
rect 49145 24395 49203 24401
rect 49145 24392 49157 24395
rect 48372 24364 49157 24392
rect 48372 24352 48378 24364
rect 49145 24361 49157 24364
rect 49191 24361 49203 24395
rect 49145 24355 49203 24361
rect 50338 24352 50344 24404
rect 50396 24392 50402 24404
rect 50801 24395 50859 24401
rect 50801 24392 50813 24395
rect 50396 24364 50813 24392
rect 50396 24352 50402 24364
rect 50801 24361 50813 24364
rect 50847 24361 50859 24395
rect 50801 24355 50859 24361
rect 36633 24327 36691 24333
rect 36633 24293 36645 24327
rect 36679 24293 36691 24327
rect 36633 24287 36691 24293
rect 36648 24256 36676 24287
rect 37366 24284 37372 24336
rect 37424 24324 37430 24336
rect 38470 24324 38476 24336
rect 37424 24296 38476 24324
rect 37424 24284 37430 24296
rect 38470 24284 38476 24296
rect 38528 24324 38534 24336
rect 38528 24296 39436 24324
rect 38528 24284 38534 24296
rect 37182 24256 37188 24268
rect 35268 24228 36676 24256
rect 37143 24228 37188 24256
rect 35268 24197 35296 24228
rect 37182 24216 37188 24228
rect 37240 24216 37246 24268
rect 38010 24256 38016 24268
rect 37923 24228 38016 24256
rect 38010 24216 38016 24228
rect 38068 24256 38074 24268
rect 39408 24256 39436 24296
rect 40034 24284 40040 24336
rect 40092 24324 40098 24336
rect 40129 24327 40187 24333
rect 40129 24324 40141 24327
rect 40092 24296 40141 24324
rect 40092 24284 40098 24296
rect 40129 24293 40141 24296
rect 40175 24324 40187 24327
rect 45370 24324 45376 24336
rect 40175 24296 45376 24324
rect 40175 24293 40187 24296
rect 40129 24287 40187 24293
rect 45370 24284 45376 24296
rect 45428 24284 45434 24336
rect 40773 24259 40831 24265
rect 40773 24256 40785 24259
rect 38068 24228 38654 24256
rect 38068 24216 38074 24228
rect 35253 24191 35311 24197
rect 35253 24157 35265 24191
rect 35299 24157 35311 24191
rect 35253 24151 35311 24157
rect 35897 24191 35955 24197
rect 35897 24157 35909 24191
rect 35943 24188 35955 24191
rect 35986 24188 35992 24200
rect 35943 24160 35992 24188
rect 35943 24157 35955 24160
rect 35897 24151 35955 24157
rect 35986 24148 35992 24160
rect 36044 24148 36050 24200
rect 37200 24188 37228 24216
rect 38197 24191 38255 24197
rect 38197 24188 38209 24191
rect 37200 24160 38209 24188
rect 38197 24157 38209 24160
rect 38243 24157 38255 24191
rect 38197 24151 38255 24157
rect 38286 24148 38292 24200
rect 38344 24188 38350 24200
rect 38626 24188 38654 24228
rect 39408 24228 40785 24256
rect 39022 24188 39028 24200
rect 38344 24160 38389 24188
rect 38626 24160 39028 24188
rect 38344 24148 38350 24160
rect 39022 24148 39028 24160
rect 39080 24148 39086 24200
rect 39408 24197 39436 24228
rect 40773 24225 40785 24228
rect 40819 24256 40831 24259
rect 40954 24256 40960 24268
rect 40819 24228 40960 24256
rect 40819 24225 40831 24228
rect 40773 24219 40831 24225
rect 40954 24216 40960 24228
rect 41012 24216 41018 24268
rect 46290 24256 46296 24268
rect 46251 24228 46296 24256
rect 46290 24216 46296 24228
rect 46348 24216 46354 24268
rect 47670 24256 47676 24268
rect 47631 24228 47676 24256
rect 47670 24216 47676 24228
rect 47728 24216 47734 24268
rect 49602 24216 49608 24268
rect 49660 24256 49666 24268
rect 50433 24259 50491 24265
rect 50433 24256 50445 24259
rect 49660 24228 50445 24256
rect 49660 24216 49666 24228
rect 50433 24225 50445 24228
rect 50479 24225 50491 24259
rect 50433 24219 50491 24225
rect 39393 24191 39451 24197
rect 39393 24157 39405 24191
rect 39439 24157 39451 24191
rect 39393 24151 39451 24157
rect 39485 24191 39543 24197
rect 39485 24157 39497 24191
rect 39531 24188 39543 24191
rect 39758 24188 39764 24200
rect 39531 24160 39764 24188
rect 39531 24157 39543 24160
rect 39485 24151 39543 24157
rect 39758 24148 39764 24160
rect 39816 24148 39822 24200
rect 39850 24148 39856 24200
rect 39908 24188 39914 24200
rect 40037 24191 40095 24197
rect 40037 24188 40049 24191
rect 39908 24160 40049 24188
rect 39908 24148 39914 24160
rect 40037 24157 40049 24160
rect 40083 24157 40095 24191
rect 40862 24188 40868 24200
rect 40775 24160 40868 24188
rect 40037 24151 40095 24157
rect 40862 24148 40868 24160
rect 40920 24148 40926 24200
rect 41509 24191 41567 24197
rect 41509 24157 41521 24191
rect 41555 24157 41567 24191
rect 41509 24151 41567 24157
rect 37001 24123 37059 24129
rect 37001 24089 37013 24123
rect 37047 24120 37059 24123
rect 37826 24120 37832 24132
rect 37047 24092 37832 24120
rect 37047 24089 37059 24092
rect 37001 24083 37059 24089
rect 37826 24080 37832 24092
rect 37884 24080 37890 24132
rect 39117 24123 39175 24129
rect 37936 24092 38884 24120
rect 35066 24052 35072 24064
rect 35027 24024 35072 24052
rect 35066 24012 35072 24024
rect 35124 24012 35130 24064
rect 37093 24055 37151 24061
rect 37093 24021 37105 24055
rect 37139 24052 37151 24055
rect 37936 24052 37964 24092
rect 38856 24064 38884 24092
rect 39117 24089 39129 24123
rect 39163 24089 39175 24123
rect 39117 24083 39175 24089
rect 39209 24123 39267 24129
rect 39209 24089 39221 24123
rect 39255 24120 39267 24123
rect 40310 24120 40316 24132
rect 39255 24092 40316 24120
rect 39255 24089 39267 24092
rect 39209 24083 39267 24089
rect 38838 24052 38844 24064
rect 37139 24024 37964 24052
rect 38799 24024 38844 24052
rect 37139 24021 37151 24024
rect 37093 24015 37151 24021
rect 38838 24012 38844 24024
rect 38896 24012 38902 24064
rect 39132 24052 39160 24083
rect 40310 24080 40316 24092
rect 40368 24120 40374 24132
rect 40880 24120 40908 24148
rect 41524 24120 41552 24151
rect 41598 24148 41604 24200
rect 41656 24188 41662 24200
rect 42705 24191 42763 24197
rect 41656 24160 41701 24188
rect 41656 24148 41662 24160
rect 42705 24157 42717 24191
rect 42751 24188 42763 24191
rect 42886 24188 42892 24200
rect 42751 24160 42892 24188
rect 42751 24157 42763 24160
rect 42705 24151 42763 24157
rect 42150 24120 42156 24132
rect 40368 24092 40908 24120
rect 41386 24092 42156 24120
rect 40368 24080 40374 24092
rect 40494 24052 40500 24064
rect 39132 24024 40500 24052
rect 40494 24012 40500 24024
rect 40552 24052 40558 24064
rect 41386 24052 41414 24092
rect 42150 24080 42156 24092
rect 42208 24120 42214 24132
rect 42720 24120 42748 24151
rect 42886 24148 42892 24160
rect 42944 24148 42950 24200
rect 43438 24148 43444 24200
rect 43496 24188 43502 24200
rect 43533 24191 43591 24197
rect 43533 24188 43545 24191
rect 43496 24160 43545 24188
rect 43496 24148 43502 24160
rect 43533 24157 43545 24160
rect 43579 24188 43591 24191
rect 45094 24188 45100 24200
rect 43579 24160 45100 24188
rect 43579 24157 43591 24160
rect 43533 24151 43591 24157
rect 45094 24148 45100 24160
rect 45152 24188 45158 24200
rect 45189 24191 45247 24197
rect 45189 24188 45201 24191
rect 45152 24160 45201 24188
rect 45152 24148 45158 24160
rect 45189 24157 45201 24160
rect 45235 24157 45247 24191
rect 45189 24151 45247 24157
rect 46569 24191 46627 24197
rect 46569 24157 46581 24191
rect 46615 24157 46627 24191
rect 47394 24188 47400 24200
rect 47355 24160 47400 24188
rect 46569 24151 46627 24157
rect 42208 24092 42748 24120
rect 44637 24123 44695 24129
rect 42208 24080 42214 24092
rect 44637 24089 44649 24123
rect 44683 24120 44695 24123
rect 46198 24120 46204 24132
rect 44683 24092 46204 24120
rect 44683 24089 44695 24092
rect 44637 24083 44695 24089
rect 46198 24080 46204 24092
rect 46256 24120 46262 24132
rect 46584 24120 46612 24151
rect 47394 24148 47400 24160
rect 47452 24148 47458 24200
rect 49694 24148 49700 24200
rect 49752 24188 49758 24200
rect 50525 24191 50583 24197
rect 50525 24188 50537 24191
rect 49752 24160 50537 24188
rect 49752 24148 49758 24160
rect 50525 24157 50537 24160
rect 50571 24157 50583 24191
rect 50525 24151 50583 24157
rect 51074 24148 51080 24200
rect 51132 24188 51138 24200
rect 51353 24191 51411 24197
rect 51353 24188 51365 24191
rect 51132 24160 51365 24188
rect 51132 24148 51138 24160
rect 51353 24157 51365 24160
rect 51399 24157 51411 24191
rect 51353 24151 51411 24157
rect 49050 24120 49056 24132
rect 46256 24092 46612 24120
rect 48898 24092 49056 24120
rect 46256 24080 46262 24092
rect 45278 24052 45284 24064
rect 40552 24024 41414 24052
rect 45239 24024 45284 24052
rect 40552 24012 40558 24024
rect 45278 24012 45284 24024
rect 45336 24012 45342 24064
rect 46290 24052 46296 24064
rect 46251 24024 46296 24052
rect 46290 24012 46296 24024
rect 46348 24012 46354 24064
rect 46584 24052 46612 24092
rect 49050 24080 49056 24092
rect 49108 24080 49114 24132
rect 49697 24055 49755 24061
rect 49697 24052 49709 24055
rect 46584 24024 49709 24052
rect 49697 24021 49709 24024
rect 49743 24052 49755 24055
rect 49878 24052 49884 24064
rect 49743 24024 49884 24052
rect 49743 24021 49755 24024
rect 49697 24015 49755 24021
rect 49878 24012 49884 24024
rect 49936 24012 49942 24064
rect 51442 24052 51448 24064
rect 51403 24024 51448 24052
rect 51442 24012 51448 24024
rect 51500 24012 51506 24064
rect 1104 23962 58880 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 58880 23962
rect 1104 23888 58880 23910
rect 34333 23851 34391 23857
rect 34333 23817 34345 23851
rect 34379 23848 34391 23851
rect 34698 23848 34704 23860
rect 34379 23820 34704 23848
rect 34379 23817 34391 23820
rect 34333 23811 34391 23817
rect 34698 23808 34704 23820
rect 34756 23808 34762 23860
rect 36538 23848 36544 23860
rect 36451 23820 36544 23848
rect 36538 23808 36544 23820
rect 36596 23848 36602 23860
rect 37182 23848 37188 23860
rect 36596 23820 37188 23848
rect 36596 23808 36602 23820
rect 37182 23808 37188 23820
rect 37240 23808 37246 23860
rect 37826 23808 37832 23860
rect 37884 23848 37890 23860
rect 37921 23851 37979 23857
rect 37921 23848 37933 23851
rect 37884 23820 37933 23848
rect 37884 23808 37890 23820
rect 37921 23817 37933 23820
rect 37967 23817 37979 23851
rect 39758 23848 39764 23860
rect 39719 23820 39764 23848
rect 37921 23811 37979 23817
rect 39758 23808 39764 23820
rect 39816 23808 39822 23860
rect 40310 23848 40316 23860
rect 40271 23820 40316 23848
rect 40310 23808 40316 23820
rect 40368 23808 40374 23860
rect 40770 23848 40776 23860
rect 40420 23820 40776 23848
rect 34716 23712 34744 23808
rect 35066 23780 35072 23792
rect 35027 23752 35072 23780
rect 35066 23740 35072 23752
rect 35124 23740 35130 23792
rect 36078 23740 36084 23792
rect 36136 23740 36142 23792
rect 38105 23783 38163 23789
rect 38105 23749 38117 23783
rect 38151 23780 38163 23783
rect 38378 23780 38384 23792
rect 38151 23752 38384 23780
rect 38151 23749 38163 23752
rect 38105 23743 38163 23749
rect 38378 23740 38384 23752
rect 38436 23780 38442 23792
rect 40420 23780 40448 23820
rect 40770 23808 40776 23820
rect 40828 23808 40834 23860
rect 41046 23808 41052 23860
rect 41104 23848 41110 23860
rect 46290 23848 46296 23860
rect 41104 23820 42748 23848
rect 41104 23808 41110 23820
rect 38436 23752 40448 23780
rect 38436 23740 38442 23752
rect 41322 23740 41328 23792
rect 41380 23740 41386 23792
rect 42720 23780 42748 23820
rect 44284 23820 46296 23848
rect 44284 23789 44312 23820
rect 46290 23808 46296 23820
rect 46348 23808 46354 23860
rect 46382 23808 46388 23860
rect 46440 23848 46446 23860
rect 47121 23851 47179 23857
rect 47121 23848 47133 23851
rect 46440 23820 47133 23848
rect 46440 23808 46446 23820
rect 47121 23817 47133 23820
rect 47167 23817 47179 23851
rect 47121 23811 47179 23817
rect 49050 23808 49056 23860
rect 49108 23848 49114 23860
rect 49145 23851 49203 23857
rect 49145 23848 49157 23851
rect 49108 23820 49157 23848
rect 49108 23808 49114 23820
rect 49145 23817 49157 23820
rect 49191 23817 49203 23851
rect 49145 23811 49203 23817
rect 44269 23783 44327 23789
rect 42720 23752 42840 23780
rect 34793 23715 34851 23721
rect 34793 23712 34805 23715
rect 34716 23684 34805 23712
rect 34793 23681 34805 23684
rect 34839 23681 34851 23715
rect 34793 23675 34851 23681
rect 37829 23715 37887 23721
rect 37829 23681 37841 23715
rect 37875 23712 37887 23715
rect 38010 23712 38016 23724
rect 37875 23684 38016 23712
rect 37875 23681 37887 23684
rect 37829 23675 37887 23681
rect 34808 23644 34836 23675
rect 38010 23672 38016 23684
rect 38068 23672 38074 23724
rect 39209 23715 39267 23721
rect 39209 23681 39221 23715
rect 39255 23712 39267 23715
rect 39850 23712 39856 23724
rect 39255 23684 39856 23712
rect 39255 23681 39267 23684
rect 39209 23675 39267 23681
rect 39850 23672 39856 23684
rect 39908 23672 39914 23724
rect 42058 23672 42064 23724
rect 42116 23712 42122 23724
rect 42702 23712 42708 23724
rect 42116 23684 42708 23712
rect 42116 23672 42122 23684
rect 42702 23672 42708 23684
rect 42760 23672 42766 23724
rect 42812 23721 42840 23752
rect 44269 23749 44281 23783
rect 44315 23749 44327 23783
rect 44269 23743 44327 23749
rect 45278 23740 45284 23792
rect 45336 23740 45342 23792
rect 46014 23780 46020 23792
rect 45975 23752 46020 23780
rect 46014 23740 46020 23752
rect 46072 23740 46078 23792
rect 49786 23780 49792 23792
rect 49747 23752 49792 23780
rect 49786 23740 49792 23752
rect 49844 23740 49850 23792
rect 51442 23780 51448 23792
rect 51106 23752 51448 23780
rect 51442 23740 51448 23752
rect 51500 23740 51506 23792
rect 42797 23715 42855 23721
rect 42797 23681 42809 23715
rect 42843 23681 42855 23715
rect 43438 23712 43444 23724
rect 43399 23684 43444 23712
rect 42797 23675 42855 23681
rect 43438 23672 43444 23684
rect 43496 23672 43502 23724
rect 46477 23715 46535 23721
rect 46477 23681 46489 23715
rect 46523 23712 46535 23715
rect 46934 23712 46940 23724
rect 46523 23684 46940 23712
rect 46523 23681 46535 23684
rect 46477 23675 46535 23681
rect 46934 23672 46940 23684
rect 46992 23672 46998 23724
rect 47762 23712 47768 23724
rect 47723 23684 47768 23712
rect 47762 23672 47768 23684
rect 47820 23672 47826 23724
rect 48041 23715 48099 23721
rect 48041 23681 48053 23715
rect 48087 23712 48099 23715
rect 48774 23712 48780 23724
rect 48087 23684 48780 23712
rect 48087 23681 48099 23684
rect 48041 23675 48099 23681
rect 48774 23672 48780 23684
rect 48832 23672 48838 23724
rect 49142 23672 49148 23724
rect 49200 23712 49206 23724
rect 49237 23715 49295 23721
rect 49237 23712 49249 23715
rect 49200 23684 49249 23712
rect 49200 23672 49206 23684
rect 49237 23681 49249 23684
rect 49283 23681 49295 23715
rect 49237 23675 49295 23681
rect 51810 23672 51816 23724
rect 51868 23712 51874 23724
rect 51868 23684 51913 23712
rect 51868 23672 51874 23684
rect 35434 23644 35440 23656
rect 34808 23616 35440 23644
rect 35434 23604 35440 23616
rect 35492 23604 35498 23656
rect 41785 23647 41843 23653
rect 41785 23613 41797 23647
rect 41831 23644 41843 23647
rect 42720 23644 42748 23672
rect 43993 23647 44051 23653
rect 43993 23644 44005 23647
rect 41831 23616 42656 23644
rect 42720 23616 44005 23644
rect 41831 23613 41843 23616
rect 41785 23607 41843 23613
rect 42628 23585 42656 23616
rect 43993 23613 44005 23616
rect 44039 23613 44051 23647
rect 43993 23607 44051 23613
rect 49878 23604 49884 23656
rect 49936 23644 49942 23656
rect 51537 23647 51595 23653
rect 51537 23644 51549 23647
rect 49936 23616 51549 23644
rect 49936 23604 49942 23616
rect 51537 23613 51549 23616
rect 51583 23613 51595 23647
rect 51537 23607 51595 23613
rect 42613 23579 42671 23585
rect 42613 23545 42625 23579
rect 42659 23545 42671 23579
rect 43349 23579 43407 23585
rect 43349 23576 43361 23579
rect 42613 23539 42671 23545
rect 42720 23548 43361 23576
rect 38105 23511 38163 23517
rect 38105 23477 38117 23511
rect 38151 23508 38163 23511
rect 38470 23508 38476 23520
rect 38151 23480 38476 23508
rect 38151 23477 38163 23480
rect 38105 23471 38163 23477
rect 38470 23468 38476 23480
rect 38528 23468 38534 23520
rect 41322 23468 41328 23520
rect 41380 23508 41386 23520
rect 42720 23508 42748 23548
rect 43349 23545 43361 23548
rect 43395 23545 43407 23579
rect 47026 23576 47032 23588
rect 43349 23539 43407 23545
rect 45296 23548 47032 23576
rect 41380 23480 42748 23508
rect 41380 23468 41386 23480
rect 42978 23468 42984 23520
rect 43036 23508 43042 23520
rect 45296 23508 45324 23548
rect 47026 23536 47032 23548
rect 47084 23536 47090 23588
rect 43036 23480 45324 23508
rect 46661 23511 46719 23517
rect 43036 23468 43042 23480
rect 46661 23477 46673 23511
rect 46707 23508 46719 23511
rect 46842 23508 46848 23520
rect 46707 23480 46848 23508
rect 46707 23477 46719 23480
rect 46661 23471 46719 23477
rect 46842 23468 46848 23480
rect 46900 23468 46906 23520
rect 49142 23468 49148 23520
rect 49200 23508 49206 23520
rect 51074 23508 51080 23520
rect 49200 23480 51080 23508
rect 49200 23468 49206 23480
rect 51074 23468 51080 23480
rect 51132 23468 51138 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 35434 23264 35440 23316
rect 35492 23304 35498 23316
rect 37829 23307 37887 23313
rect 37829 23304 37841 23307
rect 35492 23276 37841 23304
rect 35492 23264 35498 23276
rect 37829 23273 37841 23276
rect 37875 23304 37887 23307
rect 38102 23304 38108 23316
rect 37875 23276 38108 23304
rect 37875 23273 37887 23276
rect 37829 23267 37887 23273
rect 38102 23264 38108 23276
rect 38160 23264 38166 23316
rect 39117 23307 39175 23313
rect 39117 23273 39129 23307
rect 39163 23304 39175 23307
rect 41782 23304 41788 23316
rect 39163 23276 41788 23304
rect 39163 23273 39175 23276
rect 39117 23267 39175 23273
rect 41782 23264 41788 23276
rect 41840 23264 41846 23316
rect 46934 23264 46940 23316
rect 46992 23304 46998 23316
rect 47949 23307 48007 23313
rect 47949 23304 47961 23307
rect 46992 23276 47961 23304
rect 46992 23264 46998 23276
rect 47949 23273 47961 23276
rect 47995 23273 48007 23307
rect 51810 23304 51816 23316
rect 51771 23276 51816 23304
rect 47949 23267 48007 23273
rect 51810 23264 51816 23276
rect 51868 23264 51874 23316
rect 35989 23239 36047 23245
rect 35989 23205 36001 23239
rect 36035 23236 36047 23239
rect 36078 23236 36084 23248
rect 36035 23208 36084 23236
rect 36035 23205 36047 23208
rect 35989 23199 36047 23205
rect 36078 23196 36084 23208
rect 36136 23196 36142 23248
rect 44637 23239 44695 23245
rect 44637 23205 44649 23239
rect 44683 23205 44695 23239
rect 44637 23199 44695 23205
rect 49329 23239 49387 23245
rect 49329 23205 49341 23239
rect 49375 23236 49387 23239
rect 49878 23236 49884 23248
rect 49375 23208 49884 23236
rect 49375 23205 49387 23208
rect 49329 23199 49387 23205
rect 37277 23171 37335 23177
rect 37277 23137 37289 23171
rect 37323 23168 37335 23171
rect 37826 23168 37832 23180
rect 37323 23140 37832 23168
rect 37323 23137 37335 23140
rect 37277 23131 37335 23137
rect 37826 23128 37832 23140
rect 37884 23128 37890 23180
rect 39850 23168 39856 23180
rect 38672 23140 39856 23168
rect 35986 23060 35992 23112
rect 36044 23100 36050 23112
rect 36081 23103 36139 23109
rect 36081 23100 36093 23103
rect 36044 23072 36093 23100
rect 36044 23060 36050 23072
rect 36081 23069 36093 23072
rect 36127 23069 36139 23103
rect 37182 23100 37188 23112
rect 37143 23072 37188 23100
rect 36081 23063 36139 23069
rect 36096 23032 36124 23063
rect 37182 23060 37188 23072
rect 37240 23060 37246 23112
rect 37366 23100 37372 23112
rect 37327 23072 37372 23100
rect 37366 23060 37372 23072
rect 37424 23060 37430 23112
rect 38672 23109 38700 23140
rect 39850 23128 39856 23140
rect 39908 23128 39914 23180
rect 40037 23171 40095 23177
rect 40037 23137 40049 23171
rect 40083 23168 40095 23171
rect 42058 23168 42064 23180
rect 40083 23140 42064 23168
rect 40083 23137 40095 23140
rect 40037 23131 40095 23137
rect 42058 23128 42064 23140
rect 42116 23128 42122 23180
rect 38657 23103 38715 23109
rect 38657 23069 38669 23103
rect 38703 23069 38715 23103
rect 38657 23063 38715 23069
rect 38838 23060 38844 23112
rect 38896 23100 38902 23112
rect 39117 23103 39175 23109
rect 39117 23100 39129 23103
rect 38896 23072 39129 23100
rect 38896 23060 38902 23072
rect 39117 23069 39129 23072
rect 39163 23069 39175 23103
rect 39390 23100 39396 23112
rect 39351 23072 39396 23100
rect 39117 23063 39175 23069
rect 39390 23060 39396 23072
rect 39448 23060 39454 23112
rect 42978 23100 42984 23112
rect 42939 23072 42984 23100
rect 42978 23060 42984 23072
rect 43036 23060 43042 23112
rect 43809 23103 43867 23109
rect 43809 23069 43821 23103
rect 43855 23069 43867 23103
rect 43809 23063 43867 23069
rect 44453 23103 44511 23109
rect 44453 23069 44465 23103
rect 44499 23069 44511 23103
rect 44652 23100 44680 23199
rect 49878 23196 49884 23208
rect 49936 23196 49942 23248
rect 46201 23171 46259 23177
rect 46201 23137 46213 23171
rect 46247 23168 46259 23171
rect 47210 23168 47216 23180
rect 46247 23140 47216 23168
rect 46247 23137 46259 23140
rect 46201 23131 46259 23137
rect 47210 23128 47216 23140
rect 47268 23128 47274 23180
rect 48866 23168 48872 23180
rect 48827 23140 48872 23168
rect 48866 23128 48872 23140
rect 48924 23128 48930 23180
rect 45373 23103 45431 23109
rect 45373 23100 45385 23103
rect 44652 23072 45385 23100
rect 44453 23063 44511 23069
rect 45373 23069 45385 23072
rect 45419 23069 45431 23103
rect 45373 23063 45431 23069
rect 48961 23103 49019 23109
rect 48961 23069 48973 23103
rect 49007 23100 49019 23103
rect 49786 23100 49792 23112
rect 49007 23072 49792 23100
rect 49007 23069 49019 23072
rect 48961 23063 49019 23069
rect 37642 23032 37648 23044
rect 36096 23004 37648 23032
rect 37642 22992 37648 23004
rect 37700 22992 37706 23044
rect 39206 22992 39212 23044
rect 39264 23032 39270 23044
rect 40313 23035 40371 23041
rect 40313 23032 40325 23035
rect 39264 23004 40325 23032
rect 39264 22992 39270 23004
rect 40313 23001 40325 23004
rect 40359 23001 40371 23035
rect 40313 22995 40371 23001
rect 40770 22992 40776 23044
rect 40828 22992 40834 23044
rect 42061 23035 42119 23041
rect 42061 23001 42073 23035
rect 42107 23032 42119 23035
rect 42150 23032 42156 23044
rect 42107 23004 42156 23032
rect 42107 23001 42119 23004
rect 42061 22995 42119 23001
rect 42150 22992 42156 23004
rect 42208 22992 42214 23044
rect 42705 23035 42763 23041
rect 42705 23001 42717 23035
rect 42751 23032 42763 23035
rect 42794 23032 42800 23044
rect 42751 23004 42800 23032
rect 42751 23001 42763 23004
rect 42705 22995 42763 23001
rect 42794 22992 42800 23004
rect 42852 23032 42858 23044
rect 43438 23032 43444 23044
rect 42852 23004 43444 23032
rect 42852 22992 42858 23004
rect 43438 22992 43444 23004
rect 43496 23032 43502 23044
rect 43824 23032 43852 23063
rect 43496 23004 43852 23032
rect 44468 23032 44496 23063
rect 49786 23060 49792 23072
rect 49844 23060 49850 23112
rect 50246 23060 50252 23112
rect 50304 23100 50310 23112
rect 50341 23103 50399 23109
rect 50341 23100 50353 23103
rect 50304 23072 50353 23100
rect 50304 23060 50310 23072
rect 50341 23069 50353 23072
rect 50387 23069 50399 23103
rect 50341 23063 50399 23069
rect 46198 23032 46204 23044
rect 44468 23004 46204 23032
rect 43496 22992 43502 23004
rect 46198 22992 46204 23004
rect 46256 22992 46262 23044
rect 46474 23032 46480 23044
rect 46435 23004 46480 23032
rect 46474 22992 46480 23004
rect 46532 22992 46538 23044
rect 47118 22992 47124 23044
rect 47176 22992 47182 23044
rect 37274 22924 37280 22976
rect 37332 22964 37338 22976
rect 38194 22964 38200 22976
rect 37332 22936 38200 22964
rect 37332 22924 37338 22936
rect 38194 22924 38200 22936
rect 38252 22964 38258 22976
rect 38473 22967 38531 22973
rect 38473 22964 38485 22967
rect 38252 22936 38485 22964
rect 38252 22924 38258 22936
rect 38473 22933 38485 22936
rect 38519 22964 38531 22967
rect 38562 22964 38568 22976
rect 38519 22936 38568 22964
rect 38519 22933 38531 22936
rect 38473 22927 38531 22933
rect 38562 22924 38568 22936
rect 38620 22924 38626 22976
rect 39298 22964 39304 22976
rect 39259 22936 39304 22964
rect 39298 22924 39304 22936
rect 39356 22924 39362 22976
rect 43898 22964 43904 22976
rect 43859 22936 43904 22964
rect 43898 22924 43904 22936
rect 43956 22924 43962 22976
rect 44450 22924 44456 22976
rect 44508 22964 44514 22976
rect 45189 22967 45247 22973
rect 45189 22964 45201 22967
rect 44508 22936 45201 22964
rect 44508 22924 44514 22936
rect 45189 22933 45201 22936
rect 45235 22933 45247 22967
rect 45189 22927 45247 22933
rect 1104 22874 58880 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 58880 22874
rect 1104 22800 58880 22822
rect 36725 22763 36783 22769
rect 36725 22729 36737 22763
rect 36771 22729 36783 22763
rect 37550 22760 37556 22772
rect 37511 22732 37556 22760
rect 36725 22723 36783 22729
rect 36081 22627 36139 22633
rect 36081 22593 36093 22627
rect 36127 22624 36139 22627
rect 36740 22624 36768 22723
rect 37550 22720 37556 22732
rect 37608 22720 37614 22772
rect 39850 22760 39856 22772
rect 39811 22732 39856 22760
rect 39850 22720 39856 22732
rect 39908 22720 39914 22772
rect 40770 22760 40776 22772
rect 40731 22732 40776 22760
rect 40770 22720 40776 22732
rect 40828 22720 40834 22772
rect 41417 22763 41475 22769
rect 41417 22729 41429 22763
rect 41463 22760 41475 22763
rect 41506 22760 41512 22772
rect 41463 22732 41512 22760
rect 41463 22729 41475 22732
rect 41417 22723 41475 22729
rect 41506 22720 41512 22732
rect 41564 22720 41570 22772
rect 43898 22720 43904 22772
rect 43956 22760 43962 22772
rect 43956 22732 44772 22760
rect 43956 22720 43962 22732
rect 38010 22692 38016 22704
rect 37660 22664 38016 22692
rect 36127 22596 36768 22624
rect 36909 22627 36967 22633
rect 36127 22593 36139 22596
rect 36081 22587 36139 22593
rect 36909 22593 36921 22627
rect 36955 22624 36967 22627
rect 37366 22624 37372 22636
rect 36955 22596 37372 22624
rect 36955 22593 36967 22596
rect 36909 22587 36967 22593
rect 37366 22584 37372 22596
rect 37424 22584 37430 22636
rect 37660 22633 37688 22664
rect 38010 22652 38016 22664
rect 38068 22652 38074 22704
rect 39114 22652 39120 22704
rect 39172 22652 39178 22704
rect 42794 22692 42800 22704
rect 41386 22664 42800 22692
rect 37645 22627 37703 22633
rect 37645 22593 37657 22627
rect 37691 22593 37703 22627
rect 38102 22624 38108 22636
rect 38063 22596 38108 22624
rect 37645 22587 37703 22593
rect 38102 22584 38108 22596
rect 38160 22584 38166 22636
rect 40681 22627 40739 22633
rect 40681 22593 40693 22627
rect 40727 22624 40739 22627
rect 41386 22624 41414 22664
rect 42794 22652 42800 22664
rect 42852 22652 42858 22704
rect 44450 22692 44456 22704
rect 44411 22664 44456 22692
rect 44450 22652 44456 22664
rect 44508 22652 44514 22704
rect 44744 22692 44772 22732
rect 46474 22720 46480 22772
rect 46532 22760 46538 22772
rect 46661 22763 46719 22769
rect 46661 22760 46673 22763
rect 46532 22732 46673 22760
rect 46532 22720 46538 22732
rect 46661 22729 46673 22732
rect 46707 22729 46719 22763
rect 46661 22723 46719 22729
rect 49694 22720 49700 22772
rect 49752 22760 49758 22772
rect 49789 22763 49847 22769
rect 49789 22760 49801 22763
rect 49752 22732 49801 22760
rect 49752 22720 49758 22732
rect 49789 22729 49801 22732
rect 49835 22729 49847 22763
rect 49789 22723 49847 22729
rect 51074 22720 51080 22772
rect 51132 22760 51138 22772
rect 51132 22732 51177 22760
rect 51132 22720 51138 22732
rect 46198 22692 46204 22704
rect 44744 22664 44942 22692
rect 46159 22664 46204 22692
rect 46198 22652 46204 22664
rect 46256 22652 46262 22704
rect 40727 22596 41414 22624
rect 40727 22593 40739 22596
rect 40681 22587 40739 22593
rect 38378 22556 38384 22568
rect 38339 22528 38384 22556
rect 38378 22516 38384 22528
rect 38436 22516 38442 22568
rect 36262 22420 36268 22432
rect 36223 22392 36268 22420
rect 36262 22380 36268 22392
rect 36320 22380 36326 22432
rect 37642 22380 37648 22432
rect 37700 22420 37706 22432
rect 40696 22420 40724 22587
rect 42702 22584 42708 22636
rect 42760 22624 42766 22636
rect 44177 22627 44235 22633
rect 44177 22624 44189 22627
rect 42760 22596 44189 22624
rect 42760 22584 42766 22596
rect 44177 22593 44189 22596
rect 44223 22593 44235 22627
rect 46842 22624 46848 22636
rect 46803 22596 46848 22624
rect 44177 22587 44235 22593
rect 46842 22584 46848 22596
rect 46900 22584 46906 22636
rect 47394 22584 47400 22636
rect 47452 22624 47458 22636
rect 48041 22627 48099 22633
rect 48041 22624 48053 22627
rect 47452 22596 48053 22624
rect 47452 22584 47458 22596
rect 48041 22593 48053 22596
rect 48087 22593 48099 22627
rect 48041 22587 48099 22593
rect 49418 22584 49424 22636
rect 49476 22584 49482 22636
rect 50801 22627 50859 22633
rect 50801 22593 50813 22627
rect 50847 22624 50859 22627
rect 50847 22596 51074 22624
rect 50847 22593 50859 22596
rect 50801 22587 50859 22593
rect 48314 22556 48320 22568
rect 48275 22528 48320 22556
rect 48314 22516 48320 22528
rect 48372 22516 48378 22568
rect 37700 22392 40724 22420
rect 51046 22420 51074 22596
rect 51534 22420 51540 22432
rect 51046 22392 51540 22420
rect 37700 22380 37706 22392
rect 51534 22380 51540 22392
rect 51592 22420 51598 22432
rect 51721 22423 51779 22429
rect 51721 22420 51733 22423
rect 51592 22392 51733 22420
rect 51592 22380 51598 22392
rect 51721 22389 51733 22392
rect 51767 22420 51779 22423
rect 58158 22420 58164 22432
rect 51767 22392 58164 22420
rect 51767 22389 51779 22392
rect 51721 22383 51779 22389
rect 58158 22380 58164 22392
rect 58216 22380 58222 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 36262 22225 36268 22228
rect 36252 22219 36268 22225
rect 36252 22185 36264 22219
rect 36252 22179 36268 22185
rect 36262 22176 36268 22179
rect 36320 22176 36326 22228
rect 48314 22176 48320 22228
rect 48372 22216 48378 22228
rect 48501 22219 48559 22225
rect 48501 22216 48513 22219
rect 48372 22188 48513 22216
rect 48372 22176 48378 22188
rect 48501 22185 48513 22188
rect 48547 22185 48559 22219
rect 48501 22179 48559 22185
rect 37366 22108 37372 22160
rect 37424 22148 37430 22160
rect 37424 22120 38056 22148
rect 37424 22108 37430 22120
rect 35434 22080 35440 22092
rect 35395 22052 35440 22080
rect 35434 22040 35440 22052
rect 35492 22080 35498 22092
rect 38028 22089 38056 22120
rect 47780 22120 48360 22148
rect 35989 22083 36047 22089
rect 35989 22080 36001 22083
rect 35492 22052 36001 22080
rect 35492 22040 35498 22052
rect 35989 22049 36001 22052
rect 36035 22049 36047 22083
rect 35989 22043 36047 22049
rect 38013 22083 38071 22089
rect 38013 22049 38025 22083
rect 38059 22049 38071 22083
rect 38013 22043 38071 22049
rect 38565 22083 38623 22089
rect 38565 22049 38577 22083
rect 38611 22080 38623 22083
rect 39206 22080 39212 22092
rect 38611 22052 39212 22080
rect 38611 22049 38623 22052
rect 38565 22043 38623 22049
rect 39206 22040 39212 22052
rect 39264 22040 39270 22092
rect 47118 22040 47124 22092
rect 47176 22080 47182 22092
rect 47305 22083 47363 22089
rect 47305 22080 47317 22083
rect 47176 22052 47317 22080
rect 47176 22040 47182 22052
rect 47305 22049 47317 22052
rect 47351 22049 47363 22083
rect 47305 22043 47363 22049
rect 38470 22012 38476 22024
rect 38431 21984 38476 22012
rect 38470 21972 38476 21984
rect 38528 21972 38534 22024
rect 38657 22015 38715 22021
rect 38657 21981 38669 22015
rect 38703 22012 38715 22015
rect 38746 22012 38752 22024
rect 38703 21984 38752 22012
rect 38703 21981 38715 21984
rect 38657 21975 38715 21981
rect 38746 21972 38752 21984
rect 38804 21972 38810 22024
rect 39301 22015 39359 22021
rect 39301 21981 39313 22015
rect 39347 21981 39359 22015
rect 39301 21975 39359 21981
rect 37550 21944 37556 21956
rect 37490 21916 37556 21944
rect 37550 21904 37556 21916
rect 37608 21904 37614 21956
rect 38562 21904 38568 21956
rect 38620 21944 38626 21956
rect 39316 21944 39344 21975
rect 47026 21972 47032 22024
rect 47084 22012 47090 22024
rect 47213 22015 47271 22021
rect 47213 22012 47225 22015
rect 47084 21984 47225 22012
rect 47084 21972 47090 21984
rect 47213 21981 47225 21984
rect 47259 22012 47271 22015
rect 47780 22012 47808 22120
rect 48222 22080 48228 22092
rect 47872 22052 48228 22080
rect 47872 22021 47900 22052
rect 48222 22040 48228 22052
rect 48280 22040 48286 22092
rect 48332 22080 48360 22120
rect 49142 22080 49148 22092
rect 48332 22052 49148 22080
rect 49142 22040 49148 22052
rect 49200 22040 49206 22092
rect 49237 22083 49295 22089
rect 49237 22049 49249 22083
rect 49283 22080 49295 22083
rect 49418 22080 49424 22092
rect 49283 22052 49424 22080
rect 49283 22049 49295 22052
rect 49237 22043 49295 22049
rect 49418 22040 49424 22052
rect 49476 22040 49482 22092
rect 47259 21984 47808 22012
rect 47857 22015 47915 22021
rect 47259 21981 47271 21984
rect 47213 21975 47271 21981
rect 47857 21981 47869 22015
rect 47903 21981 47915 22015
rect 48685 22015 48743 22021
rect 48685 22012 48697 22015
rect 47857 21975 47915 21981
rect 48056 21984 48697 22012
rect 38620 21916 39344 21944
rect 38620 21904 38626 21916
rect 38654 21836 38660 21888
rect 38712 21876 38718 21888
rect 48056 21885 48084 21984
rect 48685 21981 48697 21984
rect 48731 21981 48743 22015
rect 49160 22012 49188 22040
rect 49329 22015 49387 22021
rect 49329 22012 49341 22015
rect 49160 21984 49341 22012
rect 48685 21975 48743 21981
rect 49329 21981 49341 21984
rect 49375 21981 49387 22015
rect 49329 21975 49387 21981
rect 39117 21879 39175 21885
rect 39117 21876 39129 21879
rect 38712 21848 39129 21876
rect 38712 21836 38718 21848
rect 39117 21845 39129 21848
rect 39163 21845 39175 21879
rect 39117 21839 39175 21845
rect 48041 21879 48099 21885
rect 48041 21845 48053 21879
rect 48087 21845 48099 21879
rect 48041 21839 48099 21845
rect 1104 21786 58880 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 58880 21786
rect 1104 21712 58880 21734
rect 37550 21672 37556 21684
rect 37511 21644 37556 21672
rect 37550 21632 37556 21644
rect 37608 21632 37614 21684
rect 38289 21675 38347 21681
rect 38289 21641 38301 21675
rect 38335 21672 38347 21675
rect 38378 21672 38384 21684
rect 38335 21644 38384 21672
rect 38335 21641 38347 21644
rect 38289 21635 38347 21641
rect 38378 21632 38384 21644
rect 38436 21632 38442 21684
rect 39114 21632 39120 21684
rect 39172 21672 39178 21684
rect 39209 21675 39267 21681
rect 39209 21672 39221 21675
rect 39172 21644 39221 21672
rect 39172 21632 39178 21644
rect 39209 21641 39221 21644
rect 39255 21641 39267 21675
rect 47762 21672 47768 21684
rect 47723 21644 47768 21672
rect 39209 21635 39267 21641
rect 47762 21632 47768 21644
rect 47820 21632 47826 21684
rect 37642 21536 37648 21548
rect 37603 21508 37648 21536
rect 37642 21496 37648 21508
rect 37700 21496 37706 21548
rect 38105 21539 38163 21545
rect 38105 21505 38117 21539
rect 38151 21536 38163 21539
rect 38654 21536 38660 21548
rect 38151 21508 38660 21536
rect 38151 21505 38163 21508
rect 38105 21499 38163 21505
rect 38654 21496 38660 21508
rect 38712 21496 38718 21548
rect 39117 21539 39175 21545
rect 39117 21505 39129 21539
rect 39163 21505 39175 21539
rect 39117 21499 39175 21505
rect 37660 21468 37688 21496
rect 39132 21468 39160 21499
rect 37660 21440 39160 21468
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 47302 21128 47308 21140
rect 47263 21100 47308 21128
rect 47302 21088 47308 21100
rect 47360 21088 47366 21140
rect 48593 20927 48651 20933
rect 48593 20893 48605 20927
rect 48639 20924 48651 20927
rect 50338 20924 50344 20936
rect 48639 20896 50344 20924
rect 48639 20893 48651 20896
rect 48593 20887 48651 20893
rect 50338 20884 50344 20896
rect 50396 20884 50402 20936
rect 1104 20698 58880 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 58880 20698
rect 1104 20624 58880 20646
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 1104 19610 58880 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 58880 19610
rect 1104 19536 58880 19558
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 1104 18522 58880 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 58880 18522
rect 1104 18448 58880 18470
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 1104 17434 58880 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 58880 17434
rect 1104 17360 58880 17382
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 1104 16346 58880 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 58880 16346
rect 1104 16272 58880 16294
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 1104 15258 58880 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 58880 15258
rect 1104 15184 58880 15206
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 1104 14170 58880 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 58880 14170
rect 1104 14096 58880 14118
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 1104 13082 58880 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 58880 13082
rect 1104 13008 58880 13030
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 1104 11994 58880 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 58880 11994
rect 1104 11920 58880 11942
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 1104 10906 58880 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 58880 10906
rect 1104 10832 58880 10854
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 1104 9818 58880 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 58880 9818
rect 1104 9744 58880 9766
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 1104 8730 58880 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 58880 8730
rect 1104 8656 58880 8678
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 1104 7642 58880 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 58880 7642
rect 1104 7568 58880 7590
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 1104 6554 58880 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 58880 6554
rect 1104 6480 58880 6502
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 1104 5466 58880 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 58880 5466
rect 1104 5392 58880 5414
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 1104 4378 58880 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 58880 4378
rect 1104 4304 58880 4326
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 1104 3290 58880 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 58880 3290
rect 1104 3216 58880 3238
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 58345 2839 58403 2845
rect 58345 2805 58357 2839
rect 58391 2836 58403 2839
rect 58618 2836 58624 2848
rect 58391 2808 58624 2836
rect 58391 2805 58403 2808
rect 58345 2799 58403 2805
rect 58618 2796 58624 2808
rect 58676 2796 58682 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 1765 2635 1823 2641
rect 1765 2601 1777 2635
rect 1811 2632 1823 2635
rect 1946 2632 1952 2644
rect 1811 2604 1952 2632
rect 1811 2601 1823 2604
rect 1765 2595 1823 2601
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 29917 2635 29975 2641
rect 29917 2601 29929 2635
rect 29963 2632 29975 2635
rect 34698 2632 34704 2644
rect 29963 2604 34704 2632
rect 29963 2601 29975 2604
rect 29917 2595 29975 2601
rect 34698 2592 34704 2604
rect 34756 2592 34762 2644
rect 58158 2632 58164 2644
rect 58119 2604 58164 2632
rect 58158 2592 58164 2604
rect 58216 2592 58222 2644
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29104 2400 29745 2428
rect 28994 2252 29000 2304
rect 29052 2292 29058 2304
rect 29104 2301 29132 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 58253 2363 58311 2369
rect 58253 2329 58265 2363
rect 58299 2360 58311 2363
rect 58618 2360 58624 2372
rect 58299 2332 58624 2360
rect 58299 2329 58311 2332
rect 58253 2323 58311 2329
rect 58618 2320 58624 2332
rect 58676 2320 58682 2372
rect 29089 2295 29147 2301
rect 29089 2292 29101 2295
rect 29052 2264 29101 2292
rect 29052 2252 29058 2264
rect 29089 2261 29101 2264
rect 29135 2261 29147 2295
rect 29089 2255 29147 2261
rect 1104 2202 58880 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 58880 2202
rect 1104 2128 58880 2150
rect 14 1300 20 1352
rect 72 1340 78 1352
rect 1578 1340 1584 1352
rect 72 1312 1584 1340
rect 72 1300 78 1312
rect 1578 1300 1584 1312
rect 1636 1300 1642 1352
<< via1 >>
rect 4874 57638 4926 57690
rect 4938 57638 4990 57690
rect 5002 57638 5054 57690
rect 5066 57638 5118 57690
rect 5130 57638 5182 57690
rect 35594 57638 35646 57690
rect 35658 57638 35710 57690
rect 35722 57638 35774 57690
rect 35786 57638 35838 57690
rect 35850 57638 35902 57690
rect 1308 57400 1360 57452
rect 1952 57196 2004 57248
rect 2044 57196 2096 57248
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 2136 56899 2188 56908
rect 2136 56865 2145 56899
rect 2145 56865 2179 56899
rect 2179 56865 2188 56899
rect 2136 56856 2188 56865
rect 1952 56831 2004 56840
rect 1952 56797 1961 56831
rect 1961 56797 1995 56831
rect 1995 56797 2004 56831
rect 1952 56788 2004 56797
rect 58348 56788 58400 56840
rect 59912 56788 59964 56840
rect 1584 56695 1636 56704
rect 1584 56661 1593 56695
rect 1593 56661 1627 56695
rect 1627 56661 1636 56695
rect 1584 56652 1636 56661
rect 2044 56695 2096 56704
rect 2044 56661 2053 56695
rect 2053 56661 2087 56695
rect 2087 56661 2096 56695
rect 2044 56652 2096 56661
rect 58624 56652 58676 56704
rect 4874 56550 4926 56602
rect 4938 56550 4990 56602
rect 5002 56550 5054 56602
rect 5066 56550 5118 56602
rect 5130 56550 5182 56602
rect 35594 56550 35646 56602
rect 35658 56550 35710 56602
rect 35722 56550 35774 56602
rect 35786 56550 35838 56602
rect 35850 56550 35902 56602
rect 30380 56448 30432 56500
rect 30932 56448 30984 56500
rect 58348 56491 58400 56500
rect 58348 56457 58357 56491
rect 58357 56457 58391 56491
rect 58391 56457 58400 56491
rect 58348 56448 58400 56457
rect 1584 56380 1636 56432
rect 2044 56108 2096 56160
rect 30380 56108 30432 56160
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 4874 55462 4926 55514
rect 4938 55462 4990 55514
rect 5002 55462 5054 55514
rect 5066 55462 5118 55514
rect 5130 55462 5182 55514
rect 35594 55462 35646 55514
rect 35658 55462 35710 55514
rect 35722 55462 35774 55514
rect 35786 55462 35838 55514
rect 35850 55462 35902 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 4874 54374 4926 54426
rect 4938 54374 4990 54426
rect 5002 54374 5054 54426
rect 5066 54374 5118 54426
rect 5130 54374 5182 54426
rect 35594 54374 35646 54426
rect 35658 54374 35710 54426
rect 35722 54374 35774 54426
rect 35786 54374 35838 54426
rect 35850 54374 35902 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 4874 53286 4926 53338
rect 4938 53286 4990 53338
rect 5002 53286 5054 53338
rect 5066 53286 5118 53338
rect 5130 53286 5182 53338
rect 35594 53286 35646 53338
rect 35658 53286 35710 53338
rect 35722 53286 35774 53338
rect 35786 53286 35838 53338
rect 35850 53286 35902 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 4874 52198 4926 52250
rect 4938 52198 4990 52250
rect 5002 52198 5054 52250
rect 5066 52198 5118 52250
rect 5130 52198 5182 52250
rect 35594 52198 35646 52250
rect 35658 52198 35710 52250
rect 35722 52198 35774 52250
rect 35786 52198 35838 52250
rect 35850 52198 35902 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 4874 51110 4926 51162
rect 4938 51110 4990 51162
rect 5002 51110 5054 51162
rect 5066 51110 5118 51162
rect 5130 51110 5182 51162
rect 35594 51110 35646 51162
rect 35658 51110 35710 51162
rect 35722 51110 35774 51162
rect 35786 51110 35838 51162
rect 35850 51110 35902 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 4874 50022 4926 50074
rect 4938 50022 4990 50074
rect 5002 50022 5054 50074
rect 5066 50022 5118 50074
rect 5130 50022 5182 50074
rect 35594 50022 35646 50074
rect 35658 50022 35710 50074
rect 35722 50022 35774 50074
rect 35786 50022 35838 50074
rect 35850 50022 35902 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 4874 48934 4926 48986
rect 4938 48934 4990 48986
rect 5002 48934 5054 48986
rect 5066 48934 5118 48986
rect 5130 48934 5182 48986
rect 35594 48934 35646 48986
rect 35658 48934 35710 48986
rect 35722 48934 35774 48986
rect 35786 48934 35838 48986
rect 35850 48934 35902 48986
rect 35348 48696 35400 48748
rect 37648 48739 37700 48748
rect 37648 48705 37657 48739
rect 37657 48705 37691 48739
rect 37691 48705 37700 48739
rect 37648 48696 37700 48705
rect 43352 48764 43404 48816
rect 40224 48696 40276 48748
rect 40592 48696 40644 48748
rect 40960 48739 41012 48748
rect 40960 48705 40969 48739
rect 40969 48705 41003 48739
rect 41003 48705 41012 48739
rect 40960 48696 41012 48705
rect 42800 48739 42852 48748
rect 42800 48705 42809 48739
rect 42809 48705 42843 48739
rect 42843 48705 42852 48739
rect 42800 48696 42852 48705
rect 36268 48671 36320 48680
rect 36268 48637 36277 48671
rect 36277 48637 36311 48671
rect 36311 48637 36320 48671
rect 36268 48628 36320 48637
rect 37556 48671 37608 48680
rect 37556 48637 37565 48671
rect 37565 48637 37599 48671
rect 37599 48637 37608 48671
rect 37556 48628 37608 48637
rect 38752 48671 38804 48680
rect 38752 48637 38761 48671
rect 38761 48637 38795 48671
rect 38795 48637 38804 48671
rect 38752 48628 38804 48637
rect 38476 48560 38528 48612
rect 43352 48560 43404 48612
rect 33140 48492 33192 48544
rect 34244 48535 34296 48544
rect 34244 48501 34253 48535
rect 34253 48501 34287 48535
rect 34287 48501 34296 48535
rect 34244 48492 34296 48501
rect 34796 48535 34848 48544
rect 34796 48501 34805 48535
rect 34805 48501 34839 48535
rect 34839 48501 34848 48535
rect 34796 48492 34848 48501
rect 38752 48492 38804 48544
rect 44272 48492 44324 48544
rect 44364 48535 44416 48544
rect 44364 48501 44373 48535
rect 44373 48501 44407 48535
rect 44407 48501 44416 48535
rect 44364 48492 44416 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 36268 48220 36320 48272
rect 37556 48220 37608 48272
rect 38476 48220 38528 48272
rect 40592 48263 40644 48272
rect 35992 48195 36044 48204
rect 32588 48084 32640 48136
rect 35992 48161 36001 48195
rect 36001 48161 36035 48195
rect 36035 48161 36044 48195
rect 35992 48152 36044 48161
rect 40132 48195 40184 48204
rect 40132 48161 40141 48195
rect 40141 48161 40175 48195
rect 40175 48161 40184 48195
rect 40132 48152 40184 48161
rect 40592 48229 40601 48263
rect 40601 48229 40635 48263
rect 40635 48229 40644 48263
rect 40592 48220 40644 48229
rect 42892 48220 42944 48272
rect 35072 48127 35124 48136
rect 35072 48093 35081 48127
rect 35081 48093 35115 48127
rect 35115 48093 35124 48127
rect 35072 48084 35124 48093
rect 34704 48016 34756 48068
rect 38752 48084 38804 48136
rect 41236 48127 41288 48136
rect 41236 48093 41245 48127
rect 41245 48093 41279 48127
rect 41279 48093 41288 48127
rect 41236 48084 41288 48093
rect 36728 48016 36780 48068
rect 33140 47991 33192 48000
rect 33140 47957 33149 47991
rect 33149 47957 33183 47991
rect 33183 47957 33192 47991
rect 33140 47948 33192 47957
rect 38292 47948 38344 48000
rect 41788 47948 41840 48000
rect 4874 47846 4926 47898
rect 4938 47846 4990 47898
rect 5002 47846 5054 47898
rect 5066 47846 5118 47898
rect 5130 47846 5182 47898
rect 35594 47846 35646 47898
rect 35658 47846 35710 47898
rect 35722 47846 35774 47898
rect 35786 47846 35838 47898
rect 35850 47846 35902 47898
rect 35072 47744 35124 47796
rect 35624 47744 35676 47796
rect 40132 47744 40184 47796
rect 33140 47676 33192 47728
rect 36084 47676 36136 47728
rect 32496 47651 32548 47660
rect 32496 47617 32505 47651
rect 32505 47617 32539 47651
rect 32539 47617 32548 47651
rect 32496 47608 32548 47617
rect 32588 47583 32640 47592
rect 32588 47549 32597 47583
rect 32597 47549 32631 47583
rect 32631 47549 32640 47583
rect 32588 47540 32640 47549
rect 31668 47472 31720 47524
rect 35532 47608 35584 47660
rect 35992 47608 36044 47660
rect 38936 47651 38988 47660
rect 38936 47617 38945 47651
rect 38945 47617 38979 47651
rect 38979 47617 38988 47651
rect 38936 47608 38988 47617
rect 37740 47583 37792 47592
rect 35348 47472 35400 47524
rect 37740 47549 37749 47583
rect 37749 47549 37783 47583
rect 37783 47549 37792 47583
rect 37740 47540 37792 47549
rect 42524 47608 42576 47660
rect 44272 47651 44324 47660
rect 44272 47617 44281 47651
rect 44281 47617 44315 47651
rect 44315 47617 44324 47651
rect 44272 47608 44324 47617
rect 44456 47651 44508 47660
rect 44456 47617 44465 47651
rect 44465 47617 44499 47651
rect 44499 47617 44508 47651
rect 44456 47608 44508 47617
rect 46480 47651 46532 47660
rect 46480 47617 46489 47651
rect 46489 47617 46523 47651
rect 46523 47617 46532 47651
rect 46480 47608 46532 47617
rect 34520 47404 34572 47456
rect 41420 47540 41472 47592
rect 42892 47583 42944 47592
rect 42892 47549 42901 47583
rect 42901 47549 42935 47583
rect 42935 47549 42944 47583
rect 42892 47540 42944 47549
rect 45836 47540 45888 47592
rect 46388 47583 46440 47592
rect 46388 47549 46397 47583
rect 46397 47549 46431 47583
rect 46431 47549 46440 47583
rect 46388 47540 46440 47549
rect 39764 47404 39816 47456
rect 41880 47447 41932 47456
rect 41880 47413 41889 47447
rect 41889 47413 41923 47447
rect 41923 47413 41932 47447
rect 41880 47404 41932 47413
rect 43076 47447 43128 47456
rect 43076 47413 43085 47447
rect 43085 47413 43119 47447
rect 43119 47413 43128 47447
rect 43076 47404 43128 47413
rect 47860 47404 47912 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 32220 47132 32272 47184
rect 38108 47200 38160 47252
rect 32864 47064 32916 47116
rect 38476 47132 38528 47184
rect 40040 47132 40092 47184
rect 41328 47132 41380 47184
rect 45008 47132 45060 47184
rect 46388 47132 46440 47184
rect 47400 47132 47452 47184
rect 37924 47064 37976 47116
rect 39856 47064 39908 47116
rect 42524 47107 42576 47116
rect 42524 47073 42533 47107
rect 42533 47073 42567 47107
rect 42567 47073 42576 47107
rect 42524 47064 42576 47073
rect 43076 47064 43128 47116
rect 45836 47064 45888 47116
rect 32220 47039 32272 47048
rect 32220 47005 32229 47039
rect 32229 47005 32263 47039
rect 32263 47005 32272 47039
rect 32220 46996 32272 47005
rect 32680 46996 32732 47048
rect 32128 46928 32180 46980
rect 32312 46860 32364 46912
rect 32956 46860 33008 46912
rect 33140 46860 33192 46912
rect 34520 46860 34572 46912
rect 35348 47039 35400 47048
rect 35348 47005 35362 47039
rect 35362 47005 35396 47039
rect 35396 47005 35400 47039
rect 35348 46996 35400 47005
rect 36176 46996 36228 47048
rect 35164 46971 35216 46980
rect 35164 46937 35173 46971
rect 35173 46937 35207 46971
rect 35207 46937 35216 46971
rect 35164 46928 35216 46937
rect 36728 46996 36780 47048
rect 37556 46996 37608 47048
rect 37464 46928 37516 46980
rect 39304 46996 39356 47048
rect 40040 47039 40092 47048
rect 40040 47005 40049 47039
rect 40049 47005 40083 47039
rect 40083 47005 40092 47039
rect 40040 46996 40092 47005
rect 38752 46928 38804 46980
rect 35624 46860 35676 46912
rect 38568 46860 38620 46912
rect 39212 46860 39264 46912
rect 40316 46903 40368 46912
rect 40316 46869 40325 46903
rect 40325 46869 40359 46903
rect 40359 46869 40368 46903
rect 40316 46860 40368 46869
rect 40408 46860 40460 46912
rect 43260 46996 43312 47048
rect 45376 47039 45428 47048
rect 45376 47005 45385 47039
rect 45385 47005 45419 47039
rect 45419 47005 45428 47039
rect 45376 46996 45428 47005
rect 41512 46860 41564 46912
rect 42984 46860 43036 46912
rect 44640 46903 44692 46912
rect 44640 46869 44649 46903
rect 44649 46869 44683 46903
rect 44683 46869 44692 46903
rect 44640 46860 44692 46869
rect 4874 46758 4926 46810
rect 4938 46758 4990 46810
rect 5002 46758 5054 46810
rect 5066 46758 5118 46810
rect 5130 46758 5182 46810
rect 35594 46758 35646 46810
rect 35658 46758 35710 46810
rect 35722 46758 35774 46810
rect 35786 46758 35838 46810
rect 35850 46758 35902 46810
rect 32588 46699 32640 46708
rect 32588 46665 32597 46699
rect 32597 46665 32631 46699
rect 32631 46665 32640 46699
rect 32588 46656 32640 46665
rect 34704 46699 34756 46708
rect 34704 46665 34713 46699
rect 34713 46665 34747 46699
rect 34747 46665 34756 46699
rect 34704 46656 34756 46665
rect 37648 46656 37700 46708
rect 38752 46656 38804 46708
rect 38936 46656 38988 46708
rect 40224 46656 40276 46708
rect 40776 46656 40828 46708
rect 31760 46520 31812 46572
rect 34244 46588 34296 46640
rect 35164 46588 35216 46640
rect 33600 46563 33652 46572
rect 33600 46529 33609 46563
rect 33609 46529 33643 46563
rect 33643 46529 33652 46563
rect 33600 46520 33652 46529
rect 34612 46563 34664 46572
rect 34612 46529 34621 46563
rect 34621 46529 34655 46563
rect 34655 46529 34664 46563
rect 34612 46520 34664 46529
rect 35532 46563 35584 46572
rect 35532 46529 35541 46563
rect 35541 46529 35575 46563
rect 35575 46529 35584 46563
rect 35532 46520 35584 46529
rect 36084 46563 36136 46572
rect 36084 46529 36093 46563
rect 36093 46529 36127 46563
rect 36127 46529 36136 46563
rect 36084 46520 36136 46529
rect 37464 46563 37516 46572
rect 37464 46529 37473 46563
rect 37473 46529 37507 46563
rect 37507 46529 37516 46563
rect 37464 46520 37516 46529
rect 37648 46563 37700 46572
rect 37648 46529 37655 46563
rect 37655 46529 37700 46563
rect 37648 46520 37700 46529
rect 40684 46588 40736 46640
rect 33324 46495 33376 46504
rect 33324 46461 33333 46495
rect 33333 46461 33367 46495
rect 33367 46461 33376 46495
rect 33324 46452 33376 46461
rect 32772 46384 32824 46436
rect 33784 46452 33836 46504
rect 37832 46563 37884 46572
rect 37832 46529 37841 46563
rect 37841 46529 37875 46563
rect 37875 46529 37884 46563
rect 37832 46520 37884 46529
rect 38016 46520 38068 46572
rect 38568 46563 38620 46572
rect 38568 46529 38577 46563
rect 38577 46529 38611 46563
rect 38611 46529 38620 46563
rect 38568 46520 38620 46529
rect 38660 46563 38712 46572
rect 38660 46529 38670 46563
rect 38670 46529 38704 46563
rect 38704 46529 38712 46563
rect 38660 46520 38712 46529
rect 39028 46563 39080 46572
rect 39028 46529 39042 46563
rect 39042 46529 39076 46563
rect 39076 46529 39080 46563
rect 39028 46520 39080 46529
rect 39212 46520 39264 46572
rect 39764 46563 39816 46572
rect 39764 46529 39774 46563
rect 39774 46529 39808 46563
rect 39808 46529 39816 46563
rect 39764 46520 39816 46529
rect 36452 46384 36504 46436
rect 37372 46384 37424 46436
rect 37832 46384 37884 46436
rect 38476 46384 38528 46436
rect 38568 46384 38620 46436
rect 40316 46520 40368 46572
rect 41420 46699 41472 46708
rect 41420 46665 41429 46699
rect 41429 46665 41463 46699
rect 41463 46665 41472 46699
rect 43260 46699 43312 46708
rect 41420 46656 41472 46665
rect 43260 46665 43269 46699
rect 43269 46665 43303 46699
rect 43303 46665 43312 46699
rect 43260 46656 43312 46665
rect 42524 46588 42576 46640
rect 42984 46631 43036 46640
rect 42984 46597 42993 46631
rect 42993 46597 43027 46631
rect 43027 46597 43036 46631
rect 42984 46588 43036 46597
rect 40224 46384 40276 46436
rect 40684 46384 40736 46436
rect 40776 46384 40828 46436
rect 42064 46520 42116 46572
rect 42708 46563 42760 46572
rect 42708 46529 42718 46563
rect 42718 46529 42752 46563
rect 42752 46529 42760 46563
rect 42708 46520 42760 46529
rect 41328 46452 41380 46504
rect 43076 46520 43128 46572
rect 43720 46588 43772 46640
rect 45376 46656 45428 46708
rect 43812 46563 43864 46572
rect 43812 46529 43821 46563
rect 43821 46529 43855 46563
rect 43855 46529 43864 46563
rect 43812 46520 43864 46529
rect 44180 46563 44232 46572
rect 43720 46452 43772 46504
rect 41512 46384 41564 46436
rect 41972 46384 42024 46436
rect 44180 46529 44189 46563
rect 44189 46529 44223 46563
rect 44223 46529 44232 46563
rect 44180 46520 44232 46529
rect 44272 46563 44324 46572
rect 44272 46529 44286 46563
rect 44286 46529 44320 46563
rect 44320 46529 44324 46563
rect 45008 46563 45060 46572
rect 44272 46520 44324 46529
rect 45008 46529 45017 46563
rect 45017 46529 45051 46563
rect 45051 46529 45060 46563
rect 45008 46520 45060 46529
rect 45100 46520 45152 46572
rect 47860 46563 47912 46572
rect 47860 46529 47869 46563
rect 47869 46529 47903 46563
rect 47903 46529 47912 46563
rect 47860 46520 47912 46529
rect 48688 46520 48740 46572
rect 48964 46520 49016 46572
rect 48780 46495 48832 46504
rect 48780 46461 48789 46495
rect 48789 46461 48823 46495
rect 48823 46461 48832 46495
rect 48780 46452 48832 46461
rect 31852 46316 31904 46368
rect 32680 46316 32732 46368
rect 33600 46316 33652 46368
rect 38660 46316 38712 46368
rect 41052 46316 41104 46368
rect 44640 46384 44692 46436
rect 48044 46384 48096 46436
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 31760 46155 31812 46164
rect 31760 46121 31769 46155
rect 31769 46121 31803 46155
rect 31803 46121 31812 46155
rect 31760 46112 31812 46121
rect 32496 46112 32548 46164
rect 34612 46112 34664 46164
rect 35532 46112 35584 46164
rect 32588 46044 32640 46096
rect 31484 45951 31536 45960
rect 31484 45917 31493 45951
rect 31493 45917 31527 45951
rect 31527 45917 31536 45951
rect 31484 45908 31536 45917
rect 32680 45976 32732 46028
rect 32128 45908 32180 45960
rect 32312 45951 32364 45960
rect 32312 45917 32321 45951
rect 32321 45917 32355 45951
rect 32355 45917 32364 45951
rect 32312 45908 32364 45917
rect 35348 46044 35400 46096
rect 33324 45976 33376 46028
rect 33416 45951 33468 45960
rect 33416 45917 33425 45951
rect 33425 45917 33459 45951
rect 33459 45917 33468 45951
rect 33416 45908 33468 45917
rect 34244 45976 34296 46028
rect 34796 45908 34848 45960
rect 34888 45908 34940 45960
rect 35900 45908 35952 45960
rect 38292 46112 38344 46164
rect 38476 46112 38528 46164
rect 40500 46112 40552 46164
rect 37648 46044 37700 46096
rect 36452 46019 36504 46028
rect 36452 45985 36461 46019
rect 36461 45985 36495 46019
rect 36495 45985 36504 46019
rect 36452 45976 36504 45985
rect 37740 46019 37792 46028
rect 37740 45985 37749 46019
rect 37749 45985 37783 46019
rect 37783 45985 37792 46019
rect 37740 45976 37792 45985
rect 38752 46044 38804 46096
rect 41236 46112 41288 46164
rect 41972 46155 42024 46164
rect 41972 46121 41981 46155
rect 41981 46121 42015 46155
rect 42015 46121 42024 46155
rect 41972 46112 42024 46121
rect 42708 46112 42760 46164
rect 43168 46112 43220 46164
rect 44180 46112 44232 46164
rect 44456 46112 44508 46164
rect 42524 46044 42576 46096
rect 43996 46044 44048 46096
rect 47032 46087 47084 46096
rect 47032 46053 47041 46087
rect 47041 46053 47075 46087
rect 47075 46053 47084 46087
rect 47032 46044 47084 46053
rect 36360 45908 36412 45960
rect 31852 45772 31904 45824
rect 32404 45772 32456 45824
rect 32956 45840 33008 45892
rect 33692 45883 33744 45892
rect 33692 45849 33701 45883
rect 33701 45849 33735 45883
rect 33735 45849 33744 45883
rect 33692 45840 33744 45849
rect 34336 45840 34388 45892
rect 36728 45951 36780 45960
rect 36728 45917 36737 45951
rect 36737 45917 36771 45951
rect 36771 45917 36780 45951
rect 36728 45908 36780 45917
rect 37556 45951 37608 45960
rect 37556 45917 37565 45951
rect 37565 45917 37599 45951
rect 37599 45917 37608 45951
rect 37556 45908 37608 45917
rect 38292 45908 38344 45960
rect 38844 45951 38896 45960
rect 38844 45917 38853 45951
rect 38853 45917 38887 45951
rect 38887 45917 38896 45951
rect 38844 45908 38896 45917
rect 40408 45951 40460 45960
rect 38660 45840 38712 45892
rect 40408 45917 40417 45951
rect 40417 45917 40451 45951
rect 40451 45917 40460 45951
rect 40408 45908 40460 45917
rect 40500 45951 40552 45960
rect 40500 45917 40510 45951
rect 40510 45917 40544 45951
rect 40544 45917 40552 45951
rect 40500 45908 40552 45917
rect 40224 45840 40276 45892
rect 43076 45976 43128 46028
rect 40868 45951 40920 45960
rect 40868 45917 40882 45951
rect 40882 45917 40916 45951
rect 40916 45917 40920 45951
rect 40868 45908 40920 45917
rect 42524 45908 42576 45960
rect 43628 45951 43680 45960
rect 43628 45917 43637 45951
rect 43637 45917 43671 45951
rect 43671 45917 43680 45951
rect 43628 45908 43680 45917
rect 44272 45908 44324 45960
rect 33048 45772 33100 45824
rect 33784 45772 33836 45824
rect 35348 45772 35400 45824
rect 38016 45772 38068 45824
rect 38752 45772 38804 45824
rect 39028 45772 39080 45824
rect 41788 45840 41840 45892
rect 44640 45840 44692 45892
rect 41972 45772 42024 45824
rect 43720 45772 43772 45824
rect 48504 45951 48556 45960
rect 48504 45917 48513 45951
rect 48513 45917 48547 45951
rect 48547 45917 48556 45951
rect 48504 45908 48556 45917
rect 48688 45951 48740 45960
rect 48688 45917 48697 45951
rect 48697 45917 48731 45951
rect 48731 45917 48740 45951
rect 48688 45908 48740 45917
rect 46204 45883 46256 45892
rect 46204 45849 46213 45883
rect 46213 45849 46247 45883
rect 46247 45849 46256 45883
rect 46204 45840 46256 45849
rect 47124 45840 47176 45892
rect 49332 45772 49384 45824
rect 49516 45815 49568 45824
rect 49516 45781 49525 45815
rect 49525 45781 49559 45815
rect 49559 45781 49568 45815
rect 49516 45772 49568 45781
rect 50804 45772 50856 45824
rect 52092 45772 52144 45824
rect 4874 45670 4926 45722
rect 4938 45670 4990 45722
rect 5002 45670 5054 45722
rect 5066 45670 5118 45722
rect 5130 45670 5182 45722
rect 35594 45670 35646 45722
rect 35658 45670 35710 45722
rect 35722 45670 35774 45722
rect 35786 45670 35838 45722
rect 35850 45670 35902 45722
rect 31852 45568 31904 45620
rect 33692 45568 33744 45620
rect 34520 45568 34572 45620
rect 36360 45568 36412 45620
rect 41972 45568 42024 45620
rect 43628 45568 43680 45620
rect 43996 45568 44048 45620
rect 48504 45568 48556 45620
rect 31576 45500 31628 45552
rect 33416 45500 33468 45552
rect 32404 45475 32456 45484
rect 32404 45441 32413 45475
rect 32413 45441 32447 45475
rect 32447 45441 32456 45475
rect 32404 45432 32456 45441
rect 33324 45475 33376 45484
rect 33324 45441 33333 45475
rect 33333 45441 33367 45475
rect 33367 45441 33376 45475
rect 33324 45432 33376 45441
rect 37648 45500 37700 45552
rect 34336 45432 34388 45484
rect 35440 45432 35492 45484
rect 36636 45475 36688 45484
rect 36636 45441 36645 45475
rect 36645 45441 36679 45475
rect 36679 45441 36688 45475
rect 36636 45432 36688 45441
rect 31852 45364 31904 45416
rect 34520 45364 34572 45416
rect 37464 45432 37516 45484
rect 37740 45432 37792 45484
rect 39212 45432 39264 45484
rect 40224 45500 40276 45552
rect 40500 45475 40552 45484
rect 40500 45441 40507 45475
rect 40507 45441 40552 45475
rect 40500 45432 40552 45441
rect 41420 45500 41472 45552
rect 34888 45296 34940 45348
rect 36176 45296 36228 45348
rect 37832 45364 37884 45416
rect 39764 45364 39816 45416
rect 37556 45296 37608 45348
rect 31116 45228 31168 45280
rect 35348 45271 35400 45280
rect 35348 45237 35357 45271
rect 35357 45237 35391 45271
rect 35391 45237 35400 45271
rect 35348 45228 35400 45237
rect 37464 45271 37516 45280
rect 37464 45237 37473 45271
rect 37473 45237 37507 45271
rect 37507 45237 37516 45271
rect 39212 45296 39264 45348
rect 40776 45475 40828 45484
rect 40776 45441 40790 45475
rect 40790 45441 40824 45475
rect 40824 45441 40828 45475
rect 40776 45432 40828 45441
rect 42800 45432 42852 45484
rect 43168 45475 43220 45484
rect 43168 45441 43177 45475
rect 43177 45441 43211 45475
rect 43211 45441 43220 45475
rect 43168 45432 43220 45441
rect 42892 45364 42944 45416
rect 47032 45500 47084 45552
rect 40960 45339 41012 45348
rect 40960 45305 40969 45339
rect 40969 45305 41003 45339
rect 41003 45305 41012 45339
rect 40960 45296 41012 45305
rect 42064 45339 42116 45348
rect 42064 45305 42073 45339
rect 42073 45305 42107 45339
rect 42107 45305 42116 45339
rect 42064 45296 42116 45305
rect 37464 45228 37516 45237
rect 38936 45228 38988 45280
rect 39304 45228 39356 45280
rect 41420 45228 41472 45280
rect 43076 45296 43128 45348
rect 45008 45475 45060 45484
rect 45008 45441 45017 45475
rect 45017 45441 45051 45475
rect 45051 45441 45060 45475
rect 45008 45432 45060 45441
rect 45100 45432 45152 45484
rect 43812 45364 43864 45416
rect 45744 45364 45796 45416
rect 49424 45432 49476 45484
rect 48412 45364 48464 45416
rect 50896 45407 50948 45416
rect 43904 45339 43956 45348
rect 42800 45228 42852 45280
rect 43904 45305 43913 45339
rect 43913 45305 43947 45339
rect 43947 45305 43956 45339
rect 43904 45296 43956 45305
rect 47952 45296 48004 45348
rect 49332 45296 49384 45348
rect 50896 45373 50905 45407
rect 50905 45373 50939 45407
rect 50939 45373 50948 45407
rect 50896 45364 50948 45373
rect 51540 45407 51592 45416
rect 51540 45373 51549 45407
rect 51549 45373 51583 45407
rect 51583 45373 51592 45407
rect 51540 45364 51592 45373
rect 50804 45296 50856 45348
rect 50528 45228 50580 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 34060 45067 34112 45076
rect 34060 45033 34069 45067
rect 34069 45033 34103 45067
rect 34103 45033 34112 45067
rect 34060 45024 34112 45033
rect 38292 45024 38344 45076
rect 31852 44931 31904 44940
rect 31852 44897 31861 44931
rect 31861 44897 31895 44931
rect 31895 44897 31904 44931
rect 31852 44888 31904 44897
rect 31116 44863 31168 44872
rect 31116 44829 31125 44863
rect 31125 44829 31159 44863
rect 31159 44829 31168 44863
rect 31116 44820 31168 44829
rect 31668 44863 31720 44872
rect 31668 44829 31677 44863
rect 31677 44829 31711 44863
rect 31711 44829 31720 44863
rect 31668 44820 31720 44829
rect 34244 44956 34296 45008
rect 34336 44956 34388 45008
rect 36084 44956 36136 45008
rect 41052 45024 41104 45076
rect 32404 44888 32456 44940
rect 34612 44888 34664 44940
rect 35348 44888 35400 44940
rect 38016 44931 38068 44940
rect 38016 44897 38025 44931
rect 38025 44897 38059 44931
rect 38059 44897 38068 44931
rect 38016 44888 38068 44897
rect 32772 44863 32824 44872
rect 32772 44829 32781 44863
rect 32781 44829 32815 44863
rect 32815 44829 32824 44863
rect 32772 44820 32824 44829
rect 32864 44820 32916 44872
rect 33508 44863 33560 44872
rect 33508 44829 33518 44863
rect 33518 44829 33552 44863
rect 33552 44829 33560 44863
rect 33508 44820 33560 44829
rect 33048 44752 33100 44804
rect 33784 44795 33836 44804
rect 33784 44761 33793 44795
rect 33793 44761 33827 44795
rect 33827 44761 33836 44795
rect 33784 44752 33836 44761
rect 32496 44684 32548 44736
rect 34520 44820 34572 44872
rect 35532 44820 35584 44872
rect 36912 44820 36964 44872
rect 37832 44863 37884 44872
rect 37832 44829 37841 44863
rect 37841 44829 37875 44863
rect 37875 44829 37884 44863
rect 37832 44820 37884 44829
rect 38292 44888 38344 44940
rect 38660 44931 38712 44940
rect 38660 44897 38669 44931
rect 38669 44897 38703 44931
rect 38703 44897 38712 44931
rect 38660 44888 38712 44897
rect 43168 45024 43220 45076
rect 43812 45067 43864 45076
rect 43812 45033 43821 45067
rect 43821 45033 43855 45067
rect 43855 45033 43864 45067
rect 43812 45024 43864 45033
rect 47124 45067 47176 45076
rect 47124 45033 47133 45067
rect 47133 45033 47167 45067
rect 47167 45033 47176 45067
rect 47124 45024 47176 45033
rect 50896 45067 50948 45076
rect 50896 45033 50905 45067
rect 50905 45033 50939 45067
rect 50939 45033 50948 45067
rect 50896 45024 50948 45033
rect 45100 44956 45152 45008
rect 43352 44931 43404 44940
rect 38200 44820 38252 44872
rect 41972 44820 42024 44872
rect 42156 44863 42208 44872
rect 42156 44829 42165 44863
rect 42165 44829 42199 44863
rect 42199 44829 42208 44863
rect 42156 44820 42208 44829
rect 42248 44863 42300 44872
rect 42248 44829 42258 44863
rect 42258 44829 42292 44863
rect 42292 44829 42300 44863
rect 42248 44820 42300 44829
rect 42432 44863 42484 44872
rect 42432 44829 42441 44863
rect 42441 44829 42475 44863
rect 42475 44829 42484 44863
rect 42432 44820 42484 44829
rect 42984 44820 43036 44872
rect 42340 44752 42392 44804
rect 43352 44897 43361 44931
rect 43361 44897 43395 44931
rect 43395 44897 43404 44931
rect 43352 44888 43404 44897
rect 49424 44888 49476 44940
rect 50620 44931 50672 44940
rect 50620 44897 50629 44931
rect 50629 44897 50663 44931
rect 50663 44897 50672 44931
rect 50620 44888 50672 44897
rect 52000 44931 52052 44940
rect 52000 44897 52009 44931
rect 52009 44897 52043 44931
rect 52043 44897 52052 44931
rect 52000 44888 52052 44897
rect 53012 44888 53064 44940
rect 43444 44863 43496 44872
rect 43444 44829 43453 44863
rect 43453 44829 43487 44863
rect 43487 44829 43496 44863
rect 43444 44820 43496 44829
rect 43996 44820 44048 44872
rect 45376 44820 45428 44872
rect 47952 44820 48004 44872
rect 50528 44863 50580 44872
rect 50528 44829 50537 44863
rect 50537 44829 50571 44863
rect 50571 44829 50580 44863
rect 50528 44820 50580 44829
rect 45008 44752 45060 44804
rect 34612 44684 34664 44736
rect 41236 44684 41288 44736
rect 42432 44684 42484 44736
rect 43628 44684 43680 44736
rect 44456 44684 44508 44736
rect 47676 44727 47728 44736
rect 47676 44693 47685 44727
rect 47685 44693 47719 44727
rect 47719 44693 47728 44727
rect 47676 44684 47728 44693
rect 49148 44684 49200 44736
rect 49240 44684 49292 44736
rect 50528 44684 50580 44736
rect 52644 44684 52696 44736
rect 4874 44582 4926 44634
rect 4938 44582 4990 44634
rect 5002 44582 5054 44634
rect 5066 44582 5118 44634
rect 5130 44582 5182 44634
rect 35594 44582 35646 44634
rect 35658 44582 35710 44634
rect 35722 44582 35774 44634
rect 35786 44582 35838 44634
rect 35850 44582 35902 44634
rect 32864 44523 32916 44532
rect 32864 44489 32873 44523
rect 32873 44489 32907 44523
rect 32907 44489 32916 44523
rect 32864 44480 32916 44489
rect 34520 44480 34572 44532
rect 38844 44480 38896 44532
rect 41420 44523 41472 44532
rect 41420 44489 41429 44523
rect 41429 44489 41463 44523
rect 41463 44489 41472 44523
rect 41420 44480 41472 44489
rect 42248 44480 42300 44532
rect 43352 44412 43404 44464
rect 43904 44480 43956 44532
rect 48412 44523 48464 44532
rect 31668 44344 31720 44396
rect 33324 44344 33376 44396
rect 34060 44344 34112 44396
rect 34520 44344 34572 44396
rect 36636 44387 36688 44396
rect 31024 44276 31076 44328
rect 32404 44276 32456 44328
rect 32956 44276 33008 44328
rect 34428 44276 34480 44328
rect 36636 44353 36645 44387
rect 36645 44353 36679 44387
rect 36679 44353 36688 44387
rect 36636 44344 36688 44353
rect 37464 44344 37516 44396
rect 38200 44387 38252 44396
rect 38200 44353 38209 44387
rect 38209 44353 38243 44387
rect 38243 44353 38252 44387
rect 38200 44344 38252 44353
rect 38936 44387 38988 44396
rect 38936 44353 38945 44387
rect 38945 44353 38979 44387
rect 38979 44353 38988 44387
rect 38936 44344 38988 44353
rect 39120 44387 39172 44396
rect 39120 44353 39129 44387
rect 39129 44353 39163 44387
rect 39163 44353 39172 44387
rect 39120 44344 39172 44353
rect 40132 44344 40184 44396
rect 37188 44276 37240 44328
rect 37740 44276 37792 44328
rect 37924 44319 37976 44328
rect 37924 44285 37933 44319
rect 37933 44285 37967 44319
rect 37967 44285 37976 44319
rect 37924 44276 37976 44285
rect 38108 44319 38160 44328
rect 38108 44285 38117 44319
rect 38117 44285 38151 44319
rect 38151 44285 38160 44319
rect 38108 44276 38160 44285
rect 40868 44276 40920 44328
rect 36912 44251 36964 44260
rect 36912 44217 36921 44251
rect 36921 44217 36955 44251
rect 36955 44217 36964 44251
rect 36912 44208 36964 44217
rect 42248 44344 42300 44396
rect 42432 44344 42484 44396
rect 42892 44387 42944 44396
rect 42892 44353 42901 44387
rect 42901 44353 42935 44387
rect 42935 44353 42944 44387
rect 42892 44344 42944 44353
rect 44456 44412 44508 44464
rect 47216 44412 47268 44464
rect 48412 44489 48421 44523
rect 48421 44489 48455 44523
rect 48455 44489 48464 44523
rect 48412 44480 48464 44489
rect 48504 44480 48556 44532
rect 49240 44480 49292 44532
rect 46940 44344 46992 44396
rect 47308 44344 47360 44396
rect 41512 44276 41564 44328
rect 43536 44319 43588 44328
rect 43536 44285 43545 44319
rect 43545 44285 43579 44319
rect 43579 44285 43588 44319
rect 43536 44276 43588 44285
rect 43996 44319 44048 44328
rect 43996 44285 44005 44319
rect 44005 44285 44039 44319
rect 44039 44285 44048 44319
rect 43996 44276 44048 44285
rect 32220 44140 32272 44192
rect 32588 44140 32640 44192
rect 36728 44140 36780 44192
rect 41236 44208 41288 44260
rect 38016 44183 38068 44192
rect 38016 44149 38025 44183
rect 38025 44149 38059 44183
rect 38059 44149 38068 44183
rect 38016 44140 38068 44149
rect 38384 44140 38436 44192
rect 39212 44140 39264 44192
rect 40684 44140 40736 44192
rect 42156 44208 42208 44260
rect 48872 44387 48924 44396
rect 48872 44353 48881 44387
rect 48881 44353 48915 44387
rect 48915 44353 48924 44387
rect 48872 44344 48924 44353
rect 48964 44387 49016 44396
rect 48964 44353 48974 44387
rect 48974 44353 49008 44387
rect 49008 44353 49016 44387
rect 49240 44387 49292 44396
rect 48964 44344 49016 44353
rect 49240 44353 49249 44387
rect 49249 44353 49283 44387
rect 49283 44353 49292 44387
rect 49240 44344 49292 44353
rect 48964 44208 49016 44260
rect 51172 44412 51224 44464
rect 50436 44387 50488 44396
rect 50436 44353 50445 44387
rect 50445 44353 50479 44387
rect 50479 44353 50488 44387
rect 50436 44344 50488 44353
rect 51724 44387 51776 44396
rect 50988 44276 51040 44328
rect 51724 44353 51733 44387
rect 51733 44353 51767 44387
rect 51767 44353 51776 44387
rect 51724 44344 51776 44353
rect 52092 44455 52144 44464
rect 52092 44421 52101 44455
rect 52101 44421 52135 44455
rect 52135 44421 52144 44455
rect 52092 44412 52144 44421
rect 51632 44276 51684 44328
rect 46296 44140 46348 44192
rect 47216 44140 47268 44192
rect 48136 44140 48188 44192
rect 50804 44208 50856 44260
rect 52828 44344 52880 44396
rect 53012 44387 53064 44396
rect 53012 44353 53021 44387
rect 53021 44353 53055 44387
rect 53055 44353 53064 44387
rect 53012 44344 53064 44353
rect 54576 44387 54628 44396
rect 52276 44208 52328 44260
rect 54576 44353 54585 44387
rect 54585 44353 54619 44387
rect 54619 44353 54628 44387
rect 54576 44344 54628 44353
rect 55772 44344 55824 44396
rect 56140 44276 56192 44328
rect 49240 44140 49292 44192
rect 50344 44140 50396 44192
rect 50528 44140 50580 44192
rect 52644 44140 52696 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 34244 43936 34296 43988
rect 36360 43936 36412 43988
rect 37096 43936 37148 43988
rect 41328 43936 41380 43988
rect 42708 43936 42760 43988
rect 43536 43936 43588 43988
rect 43812 43936 43864 43988
rect 33324 43868 33376 43920
rect 35348 43868 35400 43920
rect 36268 43868 36320 43920
rect 41144 43868 41196 43920
rect 34428 43800 34480 43852
rect 40684 43843 40736 43852
rect 31116 43732 31168 43784
rect 32680 43732 32732 43784
rect 37096 43775 37148 43784
rect 37096 43741 37105 43775
rect 37105 43741 37139 43775
rect 37139 43741 37148 43775
rect 37096 43732 37148 43741
rect 33600 43664 33652 43716
rect 34336 43664 34388 43716
rect 35072 43664 35124 43716
rect 38016 43732 38068 43784
rect 38384 43775 38436 43784
rect 38384 43741 38394 43775
rect 38394 43741 38428 43775
rect 38428 43741 38436 43775
rect 38752 43775 38804 43784
rect 38384 43732 38436 43741
rect 38752 43741 38766 43775
rect 38766 43741 38800 43775
rect 38800 43741 38804 43775
rect 38752 43732 38804 43741
rect 40684 43809 40693 43843
rect 40693 43809 40727 43843
rect 40727 43809 40736 43843
rect 40684 43800 40736 43809
rect 40592 43775 40644 43784
rect 38200 43664 38252 43716
rect 38476 43664 38528 43716
rect 33784 43596 33836 43648
rect 34060 43596 34112 43648
rect 38844 43596 38896 43648
rect 39120 43664 39172 43716
rect 40592 43741 40601 43775
rect 40601 43741 40635 43775
rect 40635 43741 40644 43775
rect 40592 43732 40644 43741
rect 41604 43800 41656 43852
rect 41328 43664 41380 43716
rect 41512 43732 41564 43784
rect 42156 43868 42208 43920
rect 45744 43911 45796 43920
rect 41972 43732 42024 43784
rect 42340 43775 42392 43784
rect 42340 43741 42347 43775
rect 42347 43741 42392 43775
rect 42340 43732 42392 43741
rect 42892 43800 42944 43852
rect 45284 43843 45336 43852
rect 45284 43809 45293 43843
rect 45293 43809 45327 43843
rect 45327 43809 45336 43843
rect 45284 43800 45336 43809
rect 45744 43877 45753 43911
rect 45753 43877 45787 43911
rect 45787 43877 45796 43911
rect 45744 43868 45796 43877
rect 46480 43936 46532 43988
rect 47032 43868 47084 43920
rect 50436 43936 50488 43988
rect 50620 43936 50672 43988
rect 51724 43936 51776 43988
rect 54576 43936 54628 43988
rect 48228 43868 48280 43920
rect 43076 43732 43128 43784
rect 45376 43775 45428 43784
rect 45376 43741 45385 43775
rect 45385 43741 45419 43775
rect 45419 43741 45428 43775
rect 45376 43732 45428 43741
rect 48964 43800 49016 43852
rect 49148 43843 49200 43852
rect 49148 43809 49157 43843
rect 49157 43809 49191 43843
rect 49191 43809 49200 43843
rect 49148 43800 49200 43809
rect 49608 43800 49660 43852
rect 50804 43868 50856 43920
rect 53932 43868 53984 43920
rect 42524 43707 42576 43716
rect 42524 43673 42533 43707
rect 42533 43673 42567 43707
rect 42567 43673 42576 43707
rect 42524 43664 42576 43673
rect 44272 43664 44324 43716
rect 47124 43707 47176 43716
rect 47124 43673 47133 43707
rect 47133 43673 47167 43707
rect 47167 43673 47176 43707
rect 47124 43664 47176 43673
rect 47216 43707 47268 43716
rect 47216 43673 47225 43707
rect 47225 43673 47259 43707
rect 47259 43673 47268 43707
rect 47492 43775 47544 43784
rect 47492 43741 47501 43775
rect 47501 43741 47535 43775
rect 47535 43741 47544 43775
rect 49240 43775 49292 43784
rect 47492 43732 47544 43741
rect 49240 43741 49249 43775
rect 49249 43741 49283 43775
rect 49283 43741 49292 43775
rect 49240 43732 49292 43741
rect 50344 43775 50396 43784
rect 50344 43741 50353 43775
rect 50353 43741 50387 43775
rect 50387 43741 50396 43775
rect 50344 43732 50396 43741
rect 50528 43775 50580 43784
rect 50528 43741 50535 43775
rect 50535 43741 50580 43775
rect 50528 43732 50580 43741
rect 51540 43800 51592 43852
rect 55496 43800 55548 43852
rect 50988 43732 51040 43784
rect 51816 43732 51868 43784
rect 53656 43775 53708 43784
rect 53656 43741 53665 43775
rect 53665 43741 53699 43775
rect 53699 43741 53708 43775
rect 53656 43732 53708 43741
rect 55312 43732 55364 43784
rect 55772 43775 55824 43784
rect 55772 43741 55781 43775
rect 55781 43741 55815 43775
rect 55815 43741 55824 43775
rect 55772 43732 55824 43741
rect 47216 43664 47268 43673
rect 39028 43596 39080 43648
rect 39396 43639 39448 43648
rect 39396 43605 39405 43639
rect 39405 43605 39439 43639
rect 39439 43605 39448 43639
rect 39396 43596 39448 43605
rect 40960 43639 41012 43648
rect 40960 43605 40969 43639
rect 40969 43605 41003 43639
rect 41003 43605 41012 43639
rect 40960 43596 41012 43605
rect 42616 43596 42668 43648
rect 42984 43596 43036 43648
rect 44180 43596 44232 43648
rect 44548 43639 44600 43648
rect 44548 43605 44557 43639
rect 44557 43605 44591 43639
rect 44591 43605 44600 43639
rect 44548 43596 44600 43605
rect 47032 43596 47084 43648
rect 47676 43664 47728 43716
rect 48780 43664 48832 43716
rect 48320 43639 48372 43648
rect 48320 43605 48329 43639
rect 48329 43605 48363 43639
rect 48363 43605 48372 43639
rect 48320 43596 48372 43605
rect 50068 43596 50120 43648
rect 50712 43707 50764 43716
rect 50712 43673 50721 43707
rect 50721 43673 50755 43707
rect 50755 43673 50764 43707
rect 50712 43664 50764 43673
rect 50896 43596 50948 43648
rect 52092 43596 52144 43648
rect 55036 43664 55088 43716
rect 53288 43596 53340 43648
rect 54484 43639 54536 43648
rect 54484 43605 54493 43639
rect 54493 43605 54527 43639
rect 54527 43605 54536 43639
rect 54484 43596 54536 43605
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 35594 43494 35646 43546
rect 35658 43494 35710 43546
rect 35722 43494 35774 43546
rect 35786 43494 35838 43546
rect 35850 43494 35902 43546
rect 34520 43392 34572 43444
rect 35348 43392 35400 43444
rect 36084 43392 36136 43444
rect 31024 43256 31076 43308
rect 32956 43299 33008 43308
rect 32956 43265 32965 43299
rect 32965 43265 32999 43299
rect 32999 43265 33008 43299
rect 32956 43256 33008 43265
rect 30012 43188 30064 43240
rect 31116 43231 31168 43240
rect 31116 43197 31125 43231
rect 31125 43197 31159 43231
rect 31159 43197 31168 43231
rect 31116 43188 31168 43197
rect 32864 43231 32916 43240
rect 32864 43197 32873 43231
rect 32873 43197 32907 43231
rect 32907 43197 32916 43231
rect 32864 43188 32916 43197
rect 33968 43299 34020 43308
rect 33968 43265 33977 43299
rect 33977 43265 34011 43299
rect 34011 43265 34020 43299
rect 33968 43256 34020 43265
rect 34796 43256 34848 43308
rect 35072 43299 35124 43308
rect 35072 43265 35082 43299
rect 35082 43265 35116 43299
rect 35116 43265 35124 43299
rect 35256 43299 35308 43308
rect 35072 43256 35124 43265
rect 35256 43265 35265 43299
rect 35265 43265 35299 43299
rect 35299 43265 35308 43299
rect 35256 43256 35308 43265
rect 36176 43324 36228 43376
rect 35532 43256 35584 43308
rect 36636 43299 36688 43308
rect 36636 43265 36645 43299
rect 36645 43265 36679 43299
rect 36679 43265 36688 43299
rect 36636 43256 36688 43265
rect 36728 43299 36780 43308
rect 36728 43265 36773 43299
rect 36773 43265 36780 43299
rect 36728 43256 36780 43265
rect 36912 43299 36964 43308
rect 36912 43265 36921 43299
rect 36921 43265 36955 43299
rect 36955 43265 36964 43299
rect 40408 43392 40460 43444
rect 40592 43435 40644 43444
rect 40592 43401 40601 43435
rect 40601 43401 40635 43435
rect 40635 43401 40644 43435
rect 40592 43392 40644 43401
rect 41604 43392 41656 43444
rect 42340 43392 42392 43444
rect 36912 43256 36964 43265
rect 34060 43188 34112 43240
rect 35624 43188 35676 43240
rect 33968 43052 34020 43104
rect 36728 43052 36780 43104
rect 37096 43052 37148 43104
rect 39304 43324 39356 43376
rect 42708 43392 42760 43444
rect 43444 43392 43496 43444
rect 46296 43435 46348 43444
rect 39212 43299 39264 43308
rect 39212 43265 39222 43299
rect 39222 43265 39256 43299
rect 39256 43265 39264 43299
rect 42524 43324 42576 43376
rect 42892 43367 42944 43376
rect 39212 43256 39264 43265
rect 40040 43299 40092 43308
rect 40040 43265 40050 43299
rect 40050 43265 40084 43299
rect 40084 43265 40092 43299
rect 40224 43299 40276 43308
rect 40040 43256 40092 43265
rect 40224 43265 40233 43299
rect 40233 43265 40267 43299
rect 40267 43265 40276 43299
rect 40224 43256 40276 43265
rect 40316 43299 40368 43308
rect 40316 43265 40325 43299
rect 40325 43265 40359 43299
rect 40359 43265 40368 43299
rect 40316 43256 40368 43265
rect 40684 43256 40736 43308
rect 41696 43299 41748 43308
rect 41696 43265 41705 43299
rect 41705 43265 41739 43299
rect 41739 43265 41748 43299
rect 41696 43256 41748 43265
rect 41788 43256 41840 43308
rect 42616 43299 42668 43308
rect 39488 43231 39540 43240
rect 39488 43197 39497 43231
rect 39497 43197 39531 43231
rect 39531 43197 39540 43231
rect 39488 43188 39540 43197
rect 39764 43188 39816 43240
rect 42616 43265 42625 43299
rect 42625 43265 42659 43299
rect 42659 43265 42668 43299
rect 42616 43256 42668 43265
rect 42892 43333 42901 43367
rect 42901 43333 42935 43367
rect 42935 43333 42944 43367
rect 42892 43324 42944 43333
rect 43628 43324 43680 43376
rect 44272 43324 44324 43376
rect 43076 43299 43128 43308
rect 43076 43265 43090 43299
rect 43090 43265 43124 43299
rect 43124 43265 43128 43299
rect 43720 43299 43772 43308
rect 43076 43256 43128 43265
rect 43720 43265 43729 43299
rect 43729 43265 43763 43299
rect 43763 43265 43772 43299
rect 43720 43256 43772 43265
rect 43904 43299 43956 43308
rect 43904 43265 43911 43299
rect 43911 43265 43956 43299
rect 43904 43256 43956 43265
rect 44180 43299 44232 43308
rect 44180 43265 44194 43299
rect 44194 43265 44228 43299
rect 44228 43265 44232 43299
rect 46296 43401 46305 43435
rect 46305 43401 46339 43435
rect 46339 43401 46348 43435
rect 46296 43392 46348 43401
rect 47492 43392 47544 43444
rect 47952 43392 48004 43444
rect 48504 43392 48556 43444
rect 52092 43392 52144 43444
rect 53932 43392 53984 43444
rect 54300 43392 54352 43444
rect 44180 43256 44232 43265
rect 38200 43120 38252 43172
rect 39304 43095 39356 43104
rect 39304 43061 39313 43095
rect 39313 43061 39347 43095
rect 39347 43061 39356 43095
rect 39304 43052 39356 43061
rect 41052 43120 41104 43172
rect 40316 43052 40368 43104
rect 44364 43188 44416 43240
rect 41972 43163 42024 43172
rect 41972 43129 41981 43163
rect 41981 43129 42015 43163
rect 42015 43129 42024 43163
rect 41972 43120 42024 43129
rect 43720 43120 43772 43172
rect 44180 43120 44232 43172
rect 41512 43052 41564 43104
rect 47032 43256 47084 43308
rect 47308 43256 47360 43308
rect 48228 43256 48280 43308
rect 48596 43256 48648 43308
rect 49608 43256 49660 43308
rect 50068 43299 50120 43308
rect 50068 43265 50077 43299
rect 50077 43265 50111 43299
rect 50111 43265 50120 43299
rect 50068 43256 50120 43265
rect 50528 43256 50580 43308
rect 51540 43299 51592 43308
rect 51540 43265 51549 43299
rect 51549 43265 51583 43299
rect 51583 43265 51592 43299
rect 51540 43256 51592 43265
rect 54944 43299 54996 43308
rect 54944 43265 54953 43299
rect 54953 43265 54987 43299
rect 54987 43265 54996 43299
rect 54944 43256 54996 43265
rect 49976 43231 50028 43240
rect 49976 43197 49985 43231
rect 49985 43197 50019 43231
rect 50019 43197 50028 43231
rect 49976 43188 50028 43197
rect 45376 43163 45428 43172
rect 45376 43129 45385 43163
rect 45385 43129 45419 43163
rect 45419 43129 45428 43163
rect 45376 43120 45428 43129
rect 46296 43120 46348 43172
rect 47952 43120 48004 43172
rect 48872 43120 48924 43172
rect 51448 43188 51500 43240
rect 55312 43231 55364 43240
rect 46940 43095 46992 43104
rect 46940 43061 46949 43095
rect 46949 43061 46983 43095
rect 46983 43061 46992 43095
rect 46940 43052 46992 43061
rect 48228 43052 48280 43104
rect 48964 43095 49016 43104
rect 48964 43061 48973 43095
rect 48973 43061 49007 43095
rect 49007 43061 49016 43095
rect 52828 43120 52880 43172
rect 55312 43197 55321 43231
rect 55321 43197 55355 43231
rect 55355 43197 55364 43231
rect 55312 43188 55364 43197
rect 55220 43120 55272 43172
rect 48964 43052 49016 43061
rect 52644 43052 52696 43104
rect 53472 43095 53524 43104
rect 53472 43061 53481 43095
rect 53481 43061 53515 43095
rect 53515 43061 53524 43095
rect 53472 43052 53524 43061
rect 55128 43052 55180 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 32956 42848 33008 42900
rect 32680 42823 32732 42832
rect 32680 42789 32689 42823
rect 32689 42789 32723 42823
rect 32723 42789 32732 42823
rect 32680 42780 32732 42789
rect 30196 42712 30248 42764
rect 31852 42712 31904 42764
rect 33324 42848 33376 42900
rect 34704 42780 34756 42832
rect 31392 42644 31444 42696
rect 31760 42644 31812 42696
rect 32220 42644 32272 42696
rect 34980 42712 35032 42764
rect 32496 42687 32548 42696
rect 32496 42653 32510 42687
rect 32510 42653 32544 42687
rect 32544 42653 32548 42687
rect 34060 42687 34112 42696
rect 32496 42644 32548 42653
rect 34060 42653 34069 42687
rect 34069 42653 34103 42687
rect 34103 42653 34112 42687
rect 34060 42644 34112 42653
rect 36452 42848 36504 42900
rect 36912 42848 36964 42900
rect 37096 42891 37148 42900
rect 37096 42857 37105 42891
rect 37105 42857 37139 42891
rect 37139 42857 37148 42891
rect 37096 42848 37148 42857
rect 36636 42780 36688 42832
rect 40224 42848 40276 42900
rect 40408 42848 40460 42900
rect 41972 42848 42024 42900
rect 42800 42848 42852 42900
rect 43444 42848 43496 42900
rect 38844 42780 38896 42832
rect 39396 42780 39448 42832
rect 43812 42780 43864 42832
rect 44640 42780 44692 42832
rect 47216 42848 47268 42900
rect 48320 42848 48372 42900
rect 48412 42848 48464 42900
rect 48872 42848 48924 42900
rect 49976 42848 50028 42900
rect 53656 42848 53708 42900
rect 54944 42848 54996 42900
rect 47124 42780 47176 42832
rect 37096 42712 37148 42764
rect 37924 42712 37976 42764
rect 39304 42712 39356 42764
rect 39672 42712 39724 42764
rect 33048 42576 33100 42628
rect 35256 42644 35308 42696
rect 35532 42687 35584 42696
rect 35532 42653 35546 42687
rect 35546 42653 35580 42687
rect 35580 42653 35584 42687
rect 35532 42644 35584 42653
rect 35992 42644 36044 42696
rect 35348 42619 35400 42628
rect 35348 42585 35357 42619
rect 35357 42585 35391 42619
rect 35391 42585 35400 42619
rect 35348 42576 35400 42585
rect 35624 42576 35676 42628
rect 34888 42508 34940 42560
rect 37832 42644 37884 42696
rect 41788 42644 41840 42696
rect 35532 42508 35584 42560
rect 36176 42508 36228 42560
rect 37188 42508 37240 42560
rect 38016 42508 38068 42560
rect 38384 42508 38436 42560
rect 40040 42551 40092 42560
rect 40040 42517 40049 42551
rect 40049 42517 40083 42551
rect 40083 42517 40092 42551
rect 40040 42508 40092 42517
rect 41696 42508 41748 42560
rect 42708 42687 42760 42696
rect 42708 42653 42717 42687
rect 42717 42653 42751 42687
rect 42751 42653 42760 42687
rect 42708 42644 42760 42653
rect 43444 42687 43496 42696
rect 43444 42653 43453 42687
rect 43453 42653 43487 42687
rect 43487 42653 43496 42687
rect 43444 42644 43496 42653
rect 44272 42712 44324 42764
rect 45008 42712 45060 42764
rect 48688 42755 48740 42764
rect 43904 42644 43956 42696
rect 44364 42644 44416 42696
rect 44548 42644 44600 42696
rect 45560 42644 45612 42696
rect 44180 42619 44232 42628
rect 44180 42585 44189 42619
rect 44189 42585 44223 42619
rect 44223 42585 44232 42619
rect 44180 42576 44232 42585
rect 44272 42576 44324 42628
rect 48688 42721 48697 42755
rect 48697 42721 48731 42755
rect 48731 42721 48740 42755
rect 48688 42712 48740 42721
rect 48044 42644 48096 42696
rect 43352 42508 43404 42560
rect 43720 42508 43772 42560
rect 48228 42576 48280 42628
rect 48872 42644 48924 42696
rect 49608 42780 49660 42832
rect 55220 42780 55272 42832
rect 51264 42712 51316 42764
rect 53380 42712 53432 42764
rect 49424 42687 49476 42696
rect 49424 42653 49433 42687
rect 49433 42653 49467 42687
rect 49467 42653 49476 42687
rect 49424 42644 49476 42653
rect 49884 42644 49936 42696
rect 52000 42687 52052 42696
rect 52000 42653 52009 42687
rect 52009 42653 52043 42687
rect 52043 42653 52052 42687
rect 52000 42644 52052 42653
rect 53104 42687 53156 42696
rect 53104 42653 53113 42687
rect 53113 42653 53147 42687
rect 53147 42653 53156 42687
rect 53104 42644 53156 42653
rect 49332 42576 49384 42628
rect 50344 42619 50396 42628
rect 50344 42585 50353 42619
rect 50353 42585 50387 42619
rect 50387 42585 50396 42619
rect 50344 42576 50396 42585
rect 53288 42644 53340 42696
rect 53472 42687 53524 42696
rect 53472 42653 53481 42687
rect 53481 42653 53515 42687
rect 53515 42653 53524 42687
rect 53472 42644 53524 42653
rect 53656 42644 53708 42696
rect 54300 42712 54352 42764
rect 54392 42687 54444 42696
rect 54392 42653 54401 42687
rect 54401 42653 54435 42687
rect 54435 42653 54444 42687
rect 54392 42644 54444 42653
rect 54760 42712 54812 42764
rect 49240 42508 49292 42560
rect 51724 42508 51776 42560
rect 53748 42576 53800 42628
rect 55128 42644 55180 42696
rect 57244 42687 57296 42696
rect 57244 42653 57253 42687
rect 57253 42653 57287 42687
rect 57287 42653 57296 42687
rect 57244 42644 57296 42653
rect 53932 42508 53984 42560
rect 54484 42508 54536 42560
rect 56692 42508 56744 42560
rect 57060 42508 57112 42560
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 35594 42406 35646 42458
rect 35658 42406 35710 42458
rect 35722 42406 35774 42458
rect 35786 42406 35838 42458
rect 35850 42406 35902 42458
rect 31760 42347 31812 42356
rect 31760 42313 31769 42347
rect 31769 42313 31803 42347
rect 31803 42313 31812 42347
rect 31760 42304 31812 42313
rect 32220 42304 32272 42356
rect 34796 42304 34848 42356
rect 34980 42304 35032 42356
rect 35992 42304 36044 42356
rect 36452 42304 36504 42356
rect 36176 42236 36228 42288
rect 38016 42304 38068 42356
rect 30012 42168 30064 42220
rect 31116 42168 31168 42220
rect 32220 42168 32272 42220
rect 34152 42168 34204 42220
rect 34612 42211 34664 42220
rect 34612 42177 34621 42211
rect 34621 42177 34655 42211
rect 34655 42177 34664 42211
rect 34612 42168 34664 42177
rect 34704 42211 34756 42220
rect 34704 42177 34713 42211
rect 34713 42177 34747 42211
rect 34747 42177 34756 42211
rect 34704 42168 34756 42177
rect 36084 42168 36136 42220
rect 38936 42211 38988 42220
rect 29276 42100 29328 42152
rect 30196 42143 30248 42152
rect 30196 42109 30205 42143
rect 30205 42109 30239 42143
rect 30239 42109 30248 42143
rect 30196 42100 30248 42109
rect 34980 42100 35032 42152
rect 35348 42100 35400 42152
rect 35440 42100 35492 42152
rect 38936 42177 38945 42211
rect 38945 42177 38979 42211
rect 38979 42177 38988 42211
rect 38936 42168 38988 42177
rect 40776 42168 40828 42220
rect 38844 42143 38896 42152
rect 38844 42109 38853 42143
rect 38853 42109 38887 42143
rect 38887 42109 38896 42143
rect 38844 42100 38896 42109
rect 32404 42032 32456 42084
rect 33692 42032 33744 42084
rect 41512 42236 41564 42288
rect 42708 42236 42760 42288
rect 41788 42211 41840 42220
rect 41788 42177 41797 42211
rect 41797 42177 41831 42211
rect 41831 42177 41840 42211
rect 41788 42168 41840 42177
rect 41880 42211 41932 42220
rect 41880 42177 41889 42211
rect 41889 42177 41923 42211
rect 41923 42177 41932 42211
rect 41880 42168 41932 42177
rect 44272 42304 44324 42356
rect 45560 42347 45612 42356
rect 45560 42313 45569 42347
rect 45569 42313 45603 42347
rect 45603 42313 45612 42347
rect 45560 42304 45612 42313
rect 47216 42304 47268 42356
rect 47860 42236 47912 42288
rect 43352 42211 43404 42220
rect 43352 42177 43361 42211
rect 43361 42177 43395 42211
rect 43395 42177 43404 42211
rect 43352 42168 43404 42177
rect 43536 42168 43588 42220
rect 43628 42211 43680 42220
rect 43628 42177 43637 42211
rect 43637 42177 43671 42211
rect 43671 42177 43680 42211
rect 43628 42168 43680 42177
rect 43904 42168 43956 42220
rect 42984 42100 43036 42152
rect 39304 42075 39356 42084
rect 39304 42041 39313 42075
rect 39313 42041 39347 42075
rect 39347 42041 39356 42075
rect 39304 42032 39356 42041
rect 32680 41964 32732 42016
rect 34152 42007 34204 42016
rect 34152 41973 34161 42007
rect 34161 41973 34195 42007
rect 34195 41973 34204 42007
rect 34152 41964 34204 41973
rect 37648 42007 37700 42016
rect 37648 41973 37657 42007
rect 37657 41973 37691 42007
rect 37691 41973 37700 42007
rect 37648 41964 37700 41973
rect 38108 41964 38160 42016
rect 38292 41964 38344 42016
rect 42340 41964 42392 42016
rect 45284 42168 45336 42220
rect 46940 42211 46992 42220
rect 46940 42177 46949 42211
rect 46949 42177 46983 42211
rect 46983 42177 46992 42211
rect 46940 42168 46992 42177
rect 47308 42168 47360 42220
rect 48964 42304 49016 42356
rect 49056 42304 49108 42356
rect 52460 42304 52512 42356
rect 52644 42304 52696 42356
rect 48136 42279 48188 42288
rect 48136 42245 48145 42279
rect 48145 42245 48179 42279
rect 48179 42245 48188 42279
rect 48136 42236 48188 42245
rect 48688 42236 48740 42288
rect 48872 42236 48924 42288
rect 48044 42211 48096 42220
rect 48044 42177 48053 42211
rect 48053 42177 48087 42211
rect 48087 42177 48096 42211
rect 48044 42168 48096 42177
rect 48228 42211 48280 42220
rect 48228 42177 48273 42211
rect 48273 42177 48280 42211
rect 48228 42168 48280 42177
rect 49240 42211 49292 42220
rect 45100 42143 45152 42152
rect 45100 42109 45109 42143
rect 45109 42109 45143 42143
rect 45143 42109 45152 42143
rect 45100 42100 45152 42109
rect 49240 42177 49249 42211
rect 49249 42177 49283 42211
rect 49283 42177 49292 42211
rect 49240 42168 49292 42177
rect 49608 42168 49660 42220
rect 49976 42168 50028 42220
rect 44272 41964 44324 42016
rect 48044 42032 48096 42084
rect 47492 41964 47544 42016
rect 48412 42032 48464 42084
rect 51080 42100 51132 42152
rect 51264 42143 51316 42152
rect 51264 42109 51273 42143
rect 51273 42109 51307 42143
rect 51307 42109 51316 42143
rect 51264 42100 51316 42109
rect 52092 42100 52144 42152
rect 53104 42304 53156 42356
rect 54760 42347 54812 42356
rect 54760 42313 54769 42347
rect 54769 42313 54803 42347
rect 54803 42313 54812 42347
rect 54760 42304 54812 42313
rect 55128 42304 55180 42356
rect 57336 42304 57388 42356
rect 53656 42236 53708 42288
rect 55036 42236 55088 42288
rect 53012 42211 53064 42220
rect 53012 42177 53021 42211
rect 53021 42177 53055 42211
rect 53055 42177 53064 42211
rect 53012 42168 53064 42177
rect 53748 42168 53800 42220
rect 54116 42211 54168 42220
rect 54116 42177 54125 42211
rect 54125 42177 54159 42211
rect 54159 42177 54168 42211
rect 54116 42168 54168 42177
rect 54300 42211 54352 42220
rect 54300 42177 54307 42211
rect 54307 42177 54352 42211
rect 54300 42168 54352 42177
rect 53196 42143 53248 42152
rect 53196 42109 53205 42143
rect 53205 42109 53239 42143
rect 53239 42109 53248 42143
rect 53196 42100 53248 42109
rect 53380 42100 53432 42152
rect 53932 42100 53984 42152
rect 54576 42211 54628 42220
rect 54576 42177 54590 42211
rect 54590 42177 54624 42211
rect 54624 42177 54628 42211
rect 54576 42168 54628 42177
rect 55036 42100 55088 42152
rect 49424 42032 49476 42084
rect 51724 42032 51776 42084
rect 49056 41964 49108 42016
rect 49700 42007 49752 42016
rect 49700 41973 49709 42007
rect 49709 41973 49743 42007
rect 49743 41973 49752 42007
rect 49700 41964 49752 41973
rect 52184 41964 52236 42016
rect 53104 41964 53156 42016
rect 54024 41964 54076 42016
rect 54392 41964 54444 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 33692 41803 33744 41812
rect 33692 41769 33701 41803
rect 33701 41769 33735 41803
rect 33735 41769 33744 41803
rect 33692 41760 33744 41769
rect 36728 41760 36780 41812
rect 40776 41803 40828 41812
rect 40776 41769 40785 41803
rect 40785 41769 40819 41803
rect 40819 41769 40828 41803
rect 40776 41760 40828 41769
rect 31024 41735 31076 41744
rect 31024 41701 31033 41735
rect 31033 41701 31067 41735
rect 31067 41701 31076 41735
rect 31024 41692 31076 41701
rect 45100 41760 45152 41812
rect 28908 41667 28960 41676
rect 28908 41633 28917 41667
rect 28917 41633 28951 41667
rect 28951 41633 28960 41667
rect 28908 41624 28960 41633
rect 30656 41624 30708 41676
rect 31852 41667 31904 41676
rect 29276 41556 29328 41608
rect 30840 41556 30892 41608
rect 31852 41633 31861 41667
rect 31861 41633 31895 41667
rect 31895 41633 31904 41667
rect 31852 41624 31904 41633
rect 33324 41667 33376 41676
rect 33324 41633 33333 41667
rect 33333 41633 33367 41667
rect 33367 41633 33376 41667
rect 33324 41624 33376 41633
rect 34704 41624 34756 41676
rect 42892 41692 42944 41744
rect 31944 41556 31996 41608
rect 32220 41599 32272 41608
rect 32220 41565 32229 41599
rect 32229 41565 32263 41599
rect 32263 41565 32272 41599
rect 32220 41556 32272 41565
rect 32772 41599 32824 41608
rect 32772 41565 32781 41599
rect 32781 41565 32815 41599
rect 32815 41565 32824 41599
rect 32772 41556 32824 41565
rect 34980 41599 35032 41608
rect 32864 41488 32916 41540
rect 34980 41565 34989 41599
rect 34989 41565 35023 41599
rect 35023 41565 35032 41599
rect 34980 41556 35032 41565
rect 37556 41624 37608 41676
rect 38016 41667 38068 41676
rect 38016 41633 38025 41667
rect 38025 41633 38059 41667
rect 38059 41633 38068 41667
rect 38016 41624 38068 41633
rect 38660 41667 38712 41676
rect 38660 41633 38669 41667
rect 38669 41633 38703 41667
rect 38703 41633 38712 41667
rect 38660 41624 38712 41633
rect 33968 41488 34020 41540
rect 37740 41556 37792 41608
rect 37924 41556 37976 41608
rect 38108 41599 38160 41608
rect 38108 41565 38117 41599
rect 38117 41565 38151 41599
rect 38151 41565 38160 41599
rect 38108 41556 38160 41565
rect 39212 41556 39264 41608
rect 40132 41599 40184 41608
rect 40132 41565 40141 41599
rect 40141 41565 40175 41599
rect 40175 41565 40184 41599
rect 40132 41556 40184 41565
rect 40224 41599 40276 41608
rect 40776 41624 40828 41676
rect 41880 41624 41932 41676
rect 40224 41565 40261 41599
rect 40261 41565 40276 41599
rect 40224 41556 40276 41565
rect 40684 41556 40736 41608
rect 40960 41556 41012 41608
rect 41328 41599 41380 41608
rect 41328 41565 41337 41599
rect 41337 41565 41371 41599
rect 41371 41565 41380 41599
rect 41328 41556 41380 41565
rect 42340 41599 42392 41608
rect 42340 41565 42349 41599
rect 42349 41565 42383 41599
rect 42383 41565 42392 41599
rect 42340 41556 42392 41565
rect 42524 41556 42576 41608
rect 43904 41667 43956 41676
rect 43904 41633 43913 41667
rect 43913 41633 43947 41667
rect 43947 41633 43956 41667
rect 43904 41624 43956 41633
rect 47584 41760 47636 41812
rect 48136 41760 48188 41812
rect 49056 41760 49108 41812
rect 49240 41760 49292 41812
rect 51080 41760 51132 41812
rect 47492 41667 47544 41676
rect 47492 41633 47501 41667
rect 47501 41633 47535 41667
rect 47535 41633 47544 41667
rect 47492 41624 47544 41633
rect 37188 41488 37240 41540
rect 40408 41531 40460 41540
rect 40408 41497 40417 41531
rect 40417 41497 40451 41531
rect 40451 41497 40460 41531
rect 40408 41488 40460 41497
rect 37648 41420 37700 41472
rect 42248 41488 42300 41540
rect 47400 41599 47452 41608
rect 47400 41565 47409 41599
rect 47409 41565 47443 41599
rect 47443 41565 47452 41599
rect 47400 41556 47452 41565
rect 48320 41599 48372 41608
rect 48320 41565 48329 41599
rect 48329 41565 48363 41599
rect 48363 41565 48372 41599
rect 48320 41556 48372 41565
rect 49056 41556 49108 41608
rect 51908 41692 51960 41744
rect 52092 41692 52144 41744
rect 49700 41624 49752 41676
rect 51540 41624 51592 41676
rect 50528 41599 50580 41608
rect 50528 41565 50537 41599
rect 50537 41565 50571 41599
rect 50571 41565 50580 41599
rect 50528 41556 50580 41565
rect 51172 41556 51224 41608
rect 52184 41599 52236 41608
rect 52184 41565 52194 41599
rect 52194 41565 52228 41599
rect 52228 41565 52236 41599
rect 52644 41624 52696 41676
rect 52184 41556 52236 41565
rect 52828 41556 52880 41608
rect 53104 41624 53156 41676
rect 53564 41624 53616 41676
rect 54024 41667 54076 41676
rect 54024 41633 54033 41667
rect 54033 41633 54067 41667
rect 54067 41633 54076 41667
rect 54024 41624 54076 41633
rect 57244 41624 57296 41676
rect 57428 41624 57480 41676
rect 53932 41599 53984 41608
rect 53932 41565 53941 41599
rect 53941 41565 53975 41599
rect 53975 41565 53984 41599
rect 53932 41556 53984 41565
rect 56232 41599 56284 41608
rect 43076 41488 43128 41540
rect 48780 41488 48832 41540
rect 49240 41488 49292 41540
rect 43720 41420 43772 41472
rect 47952 41420 48004 41472
rect 49608 41488 49660 41540
rect 49792 41420 49844 41472
rect 49976 41420 50028 41472
rect 50896 41463 50948 41472
rect 50896 41429 50905 41463
rect 50905 41429 50939 41463
rect 50939 41429 50948 41463
rect 50896 41420 50948 41429
rect 50988 41420 51040 41472
rect 51724 41420 51776 41472
rect 52000 41420 52052 41472
rect 52276 41488 52328 41540
rect 56232 41565 56241 41599
rect 56241 41565 56275 41599
rect 56275 41565 56284 41599
rect 56232 41556 56284 41565
rect 53840 41420 53892 41472
rect 54392 41488 54444 41540
rect 54300 41420 54352 41472
rect 54484 41420 54536 41472
rect 55036 41420 55088 41472
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 35594 41318 35646 41370
rect 35658 41318 35710 41370
rect 35722 41318 35774 41370
rect 35786 41318 35838 41370
rect 35850 41318 35902 41370
rect 32312 41080 32364 41132
rect 34980 41216 35032 41268
rect 36636 41216 36688 41268
rect 37464 41216 37516 41268
rect 34796 41148 34848 41200
rect 38384 41216 38436 41268
rect 33324 41080 33376 41132
rect 35440 41123 35492 41132
rect 35440 41089 35444 41123
rect 35444 41089 35478 41123
rect 35478 41089 35492 41123
rect 35440 41080 35492 41089
rect 35532 41123 35584 41132
rect 35532 41089 35541 41123
rect 35541 41089 35575 41123
rect 35575 41089 35584 41123
rect 35808 41123 35860 41132
rect 35532 41080 35584 41089
rect 35808 41089 35816 41123
rect 35816 41089 35850 41123
rect 35850 41089 35860 41123
rect 35808 41080 35860 41089
rect 35900 41123 35952 41132
rect 35900 41089 35909 41123
rect 35909 41089 35943 41123
rect 35943 41089 35952 41123
rect 35900 41080 35952 41089
rect 37280 41080 37332 41132
rect 37556 41123 37608 41132
rect 37556 41089 37565 41123
rect 37565 41089 37599 41123
rect 37599 41089 37608 41123
rect 37556 41080 37608 41089
rect 38108 41148 38160 41200
rect 38568 41216 38620 41268
rect 38936 41216 38988 41268
rect 44272 41216 44324 41268
rect 47860 41259 47912 41268
rect 47860 41225 47869 41259
rect 47869 41225 47903 41259
rect 47903 41225 47912 41259
rect 47860 41216 47912 41225
rect 48228 41216 48280 41268
rect 49240 41259 49292 41268
rect 49240 41225 49249 41259
rect 49249 41225 49283 41259
rect 49283 41225 49292 41259
rect 49240 41216 49292 41225
rect 50252 41216 50304 41268
rect 51080 41216 51132 41268
rect 37924 41080 37976 41132
rect 38384 41080 38436 41132
rect 38614 41123 38666 41132
rect 38614 41089 38640 41123
rect 38640 41089 38666 41123
rect 38614 41080 38666 41089
rect 38752 41080 38804 41132
rect 29092 41012 29144 41064
rect 40684 41080 40736 41132
rect 35440 40944 35492 40996
rect 35992 40944 36044 40996
rect 37740 40987 37792 40996
rect 37740 40953 37749 40987
rect 37749 40953 37783 40987
rect 37783 40953 37792 40987
rect 37740 40944 37792 40953
rect 38568 40944 38620 40996
rect 39488 40944 39540 40996
rect 40776 40944 40828 40996
rect 42340 41148 42392 41200
rect 42524 41148 42576 41200
rect 43996 41148 44048 41200
rect 41696 41080 41748 41132
rect 41972 41080 42024 41132
rect 42340 40944 42392 40996
rect 43168 41080 43220 41132
rect 43904 41123 43956 41132
rect 43904 41089 43913 41123
rect 43913 41089 43947 41123
rect 43947 41089 43956 41123
rect 43904 41080 43956 41089
rect 46664 41080 46716 41132
rect 48320 41080 48372 41132
rect 42984 41012 43036 41064
rect 36636 40876 36688 40928
rect 37556 40876 37608 40928
rect 38108 40876 38160 40928
rect 39672 40876 39724 40928
rect 40132 40876 40184 40928
rect 42248 40876 42300 40928
rect 48872 41012 48924 41064
rect 49332 41080 49384 41132
rect 49608 41080 49660 41132
rect 50252 41055 50304 41064
rect 50252 41021 50261 41055
rect 50261 41021 50295 41055
rect 50295 41021 50304 41055
rect 50252 41012 50304 41021
rect 48412 40944 48464 40996
rect 49608 40944 49660 40996
rect 51724 41191 51776 41200
rect 51724 41157 51733 41191
rect 51733 41157 51767 41191
rect 51767 41157 51776 41191
rect 51724 41148 51776 41157
rect 51908 41148 51960 41200
rect 54392 41148 54444 41200
rect 54760 41148 54812 41200
rect 50804 41123 50856 41132
rect 50804 41089 50813 41123
rect 50813 41089 50847 41123
rect 50847 41089 50856 41123
rect 50804 41080 50856 41089
rect 51632 41080 51684 41132
rect 51816 41123 51868 41132
rect 51816 41089 51821 41123
rect 51821 41089 51855 41123
rect 51855 41089 51868 41123
rect 51816 41080 51868 41089
rect 52000 41080 52052 41132
rect 52368 41080 52420 41132
rect 53840 41123 53892 41132
rect 53840 41089 53849 41123
rect 53849 41089 53883 41123
rect 53883 41089 53892 41123
rect 53840 41080 53892 41089
rect 54024 41080 54076 41132
rect 56232 41216 56284 41268
rect 54484 41012 54536 41064
rect 54668 41012 54720 41064
rect 55588 41012 55640 41064
rect 54576 40944 54628 40996
rect 48964 40876 49016 40928
rect 51172 40876 51224 40928
rect 52000 40876 52052 40928
rect 53104 40919 53156 40928
rect 53104 40885 53113 40919
rect 53113 40885 53147 40919
rect 53147 40885 53156 40919
rect 53104 40876 53156 40885
rect 53932 40876 53984 40928
rect 55036 40876 55088 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 29092 40715 29144 40724
rect 29092 40681 29101 40715
rect 29101 40681 29135 40715
rect 29135 40681 29144 40715
rect 29092 40672 29144 40681
rect 30840 40672 30892 40724
rect 32404 40672 32456 40724
rect 34704 40672 34756 40724
rect 35900 40672 35952 40724
rect 36636 40672 36688 40724
rect 36728 40672 36780 40724
rect 37924 40715 37976 40724
rect 37924 40681 37933 40715
rect 37933 40681 37967 40715
rect 37967 40681 37976 40715
rect 37924 40672 37976 40681
rect 38476 40672 38528 40724
rect 40040 40672 40092 40724
rect 45008 40672 45060 40724
rect 29828 40536 29880 40588
rect 28908 40468 28960 40520
rect 30564 40511 30616 40520
rect 30564 40477 30573 40511
rect 30573 40477 30607 40511
rect 30607 40477 30616 40511
rect 30564 40468 30616 40477
rect 32404 40536 32456 40588
rect 30380 40400 30432 40452
rect 31760 40468 31812 40520
rect 32772 40468 32824 40520
rect 30840 40443 30892 40452
rect 30840 40409 30849 40443
rect 30849 40409 30883 40443
rect 30883 40409 30892 40443
rect 30840 40400 30892 40409
rect 30932 40443 30984 40452
rect 30932 40409 30941 40443
rect 30941 40409 30975 40443
rect 30975 40409 30984 40443
rect 30932 40400 30984 40409
rect 31852 40400 31904 40452
rect 32588 40400 32640 40452
rect 33232 40511 33284 40520
rect 33232 40477 33241 40511
rect 33241 40477 33275 40511
rect 33275 40477 33284 40511
rect 35532 40604 35584 40656
rect 40776 40604 40828 40656
rect 42708 40604 42760 40656
rect 35348 40579 35400 40588
rect 35348 40545 35357 40579
rect 35357 40545 35391 40579
rect 35391 40545 35400 40579
rect 35348 40536 35400 40545
rect 33232 40468 33284 40477
rect 35256 40468 35308 40520
rect 37188 40536 37240 40588
rect 37832 40579 37884 40588
rect 37832 40545 37841 40579
rect 37841 40545 37875 40579
rect 37875 40545 37884 40579
rect 37832 40536 37884 40545
rect 54116 40672 54168 40724
rect 45284 40579 45336 40588
rect 36728 40468 36780 40520
rect 37004 40468 37056 40520
rect 39212 40468 39264 40520
rect 40684 40511 40736 40520
rect 40684 40477 40693 40511
rect 40693 40477 40727 40511
rect 40727 40477 40736 40511
rect 40684 40468 40736 40477
rect 37648 40400 37700 40452
rect 37924 40400 37976 40452
rect 32956 40375 33008 40384
rect 32956 40341 32965 40375
rect 32965 40341 32999 40375
rect 32999 40341 33008 40375
rect 32956 40332 33008 40341
rect 37096 40375 37148 40384
rect 37096 40341 37105 40375
rect 37105 40341 37139 40375
rect 37139 40341 37148 40375
rect 37096 40332 37148 40341
rect 37188 40332 37240 40384
rect 39488 40400 39540 40452
rect 40040 40332 40092 40384
rect 40500 40332 40552 40384
rect 45284 40545 45293 40579
rect 45293 40545 45327 40579
rect 45327 40545 45336 40579
rect 45284 40536 45336 40545
rect 48136 40604 48188 40656
rect 48412 40604 48464 40656
rect 51540 40604 51592 40656
rect 48320 40536 48372 40588
rect 50896 40579 50948 40588
rect 41696 40468 41748 40520
rect 45468 40468 45520 40520
rect 46664 40511 46716 40520
rect 46664 40477 46673 40511
rect 46673 40477 46707 40511
rect 46707 40477 46716 40511
rect 46664 40468 46716 40477
rect 50896 40545 50905 40579
rect 50905 40545 50939 40579
rect 50939 40545 50948 40579
rect 50896 40536 50948 40545
rect 51172 40536 51224 40588
rect 41972 40400 42024 40452
rect 45192 40400 45244 40452
rect 42064 40332 42116 40384
rect 47492 40375 47544 40384
rect 47492 40341 47501 40375
rect 47501 40341 47535 40375
rect 47535 40341 47544 40375
rect 47492 40332 47544 40341
rect 48320 40375 48372 40384
rect 48320 40341 48329 40375
rect 48329 40341 48363 40375
rect 48363 40341 48372 40375
rect 48320 40332 48372 40341
rect 48780 40511 48832 40520
rect 48780 40477 48825 40511
rect 48825 40477 48832 40511
rect 48780 40468 48832 40477
rect 48964 40511 49016 40520
rect 48964 40477 48973 40511
rect 48973 40477 49007 40511
rect 49007 40477 49016 40511
rect 48964 40468 49016 40477
rect 49516 40468 49568 40520
rect 52000 40511 52052 40520
rect 52000 40477 52009 40511
rect 52009 40477 52043 40511
rect 52043 40477 52052 40511
rect 52000 40468 52052 40477
rect 52092 40511 52144 40520
rect 52092 40477 52102 40511
rect 52102 40477 52136 40511
rect 52136 40477 52144 40511
rect 52368 40511 52420 40520
rect 52092 40468 52144 40477
rect 52368 40477 52377 40511
rect 52377 40477 52411 40511
rect 52411 40477 52420 40511
rect 52368 40468 52420 40477
rect 53656 40536 53708 40588
rect 53840 40536 53892 40588
rect 49424 40400 49476 40452
rect 49884 40400 49936 40452
rect 51264 40400 51316 40452
rect 52276 40443 52328 40452
rect 49700 40375 49752 40384
rect 49700 40341 49709 40375
rect 49709 40341 49743 40375
rect 49743 40341 49752 40375
rect 49700 40332 49752 40341
rect 51172 40332 51224 40384
rect 51448 40375 51500 40384
rect 51448 40341 51457 40375
rect 51457 40341 51491 40375
rect 51491 40341 51500 40375
rect 51448 40332 51500 40341
rect 52276 40409 52285 40443
rect 52285 40409 52319 40443
rect 52319 40409 52328 40443
rect 52276 40400 52328 40409
rect 52828 40400 52880 40452
rect 53380 40468 53432 40520
rect 53932 40511 53984 40520
rect 53932 40477 53941 40511
rect 53941 40477 53975 40511
rect 53975 40477 53984 40511
rect 53932 40468 53984 40477
rect 54024 40511 54076 40520
rect 54024 40477 54034 40511
rect 54034 40477 54068 40511
rect 54068 40477 54076 40511
rect 54300 40536 54352 40588
rect 54024 40468 54076 40477
rect 54576 40468 54628 40520
rect 55588 40511 55640 40520
rect 55588 40477 55597 40511
rect 55597 40477 55631 40511
rect 55631 40477 55640 40511
rect 55588 40468 55640 40477
rect 57244 40511 57296 40520
rect 57244 40477 57253 40511
rect 57253 40477 57287 40511
rect 57287 40477 57296 40511
rect 57244 40468 57296 40477
rect 57428 40511 57480 40520
rect 57428 40477 57437 40511
rect 57437 40477 57471 40511
rect 57471 40477 57480 40511
rect 57428 40468 57480 40477
rect 54484 40400 54536 40452
rect 55036 40400 55088 40452
rect 56600 40443 56652 40452
rect 56600 40409 56609 40443
rect 56609 40409 56643 40443
rect 56643 40409 56652 40443
rect 56600 40400 56652 40409
rect 53104 40332 53156 40384
rect 54852 40332 54904 40384
rect 58256 40375 58308 40384
rect 58256 40341 58265 40375
rect 58265 40341 58299 40375
rect 58299 40341 58308 40375
rect 58256 40332 58308 40341
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 35594 40230 35646 40282
rect 35658 40230 35710 40282
rect 35722 40230 35774 40282
rect 35786 40230 35838 40282
rect 35850 40230 35902 40282
rect 30840 40128 30892 40180
rect 31576 40128 31628 40180
rect 30656 39992 30708 40044
rect 30932 40035 30984 40044
rect 30932 40001 30939 40035
rect 30939 40001 30984 40035
rect 30932 39992 30984 40001
rect 31116 40035 31168 40044
rect 31116 40001 31125 40035
rect 31125 40001 31159 40035
rect 31159 40001 31168 40035
rect 31116 39992 31168 40001
rect 31760 40060 31812 40112
rect 38108 40128 38160 40180
rect 40408 40128 40460 40180
rect 32496 40035 32548 40044
rect 29184 39924 29236 39976
rect 30380 39924 30432 39976
rect 32496 40001 32500 40035
rect 32500 40001 32534 40035
rect 32534 40001 32548 40035
rect 32496 39992 32548 40001
rect 33232 40060 33284 40112
rect 34612 40060 34664 40112
rect 37740 40103 37792 40112
rect 37740 40069 37749 40103
rect 37749 40069 37783 40103
rect 37783 40069 37792 40103
rect 37740 40060 37792 40069
rect 32956 40035 33008 40044
rect 32956 40001 32965 40035
rect 32965 40001 32999 40035
rect 32999 40001 33008 40035
rect 33600 40035 33652 40044
rect 32956 39992 33008 40001
rect 33600 40001 33609 40035
rect 33609 40001 33643 40035
rect 33643 40001 33652 40035
rect 33600 39992 33652 40001
rect 36084 40035 36136 40044
rect 36084 40001 36093 40035
rect 36093 40001 36127 40035
rect 36127 40001 36136 40035
rect 36084 39992 36136 40001
rect 37096 39992 37148 40044
rect 37648 40035 37700 40044
rect 37648 40001 37655 40035
rect 37655 40001 37700 40035
rect 37648 39992 37700 40001
rect 33508 39967 33560 39976
rect 33508 39933 33517 39967
rect 33517 39933 33551 39967
rect 33551 39933 33560 39967
rect 33508 39924 33560 39933
rect 34060 39924 34112 39976
rect 31392 39899 31444 39908
rect 31392 39865 31401 39899
rect 31401 39865 31435 39899
rect 31435 39865 31444 39899
rect 31392 39856 31444 39865
rect 32312 39899 32364 39908
rect 32312 39865 32321 39899
rect 32321 39865 32355 39899
rect 32355 39865 32364 39899
rect 32312 39856 32364 39865
rect 33968 39899 34020 39908
rect 33968 39865 33977 39899
rect 33977 39865 34011 39899
rect 34011 39865 34020 39899
rect 33968 39856 34020 39865
rect 29000 39788 29052 39840
rect 32220 39788 32272 39840
rect 35256 39788 35308 39840
rect 35532 39788 35584 39840
rect 36912 39856 36964 39908
rect 37924 39992 37976 40044
rect 38568 39992 38620 40044
rect 38108 39924 38160 39976
rect 41972 40103 42024 40112
rect 38844 39992 38896 40044
rect 39856 40035 39908 40044
rect 39856 40001 39865 40035
rect 39865 40001 39899 40035
rect 39899 40001 39908 40035
rect 39856 39992 39908 40001
rect 41696 40035 41748 40044
rect 41696 40001 41705 40035
rect 41705 40001 41739 40035
rect 41739 40001 41748 40035
rect 41696 39992 41748 40001
rect 41972 40069 41981 40103
rect 41981 40069 42015 40103
rect 42015 40069 42024 40103
rect 41972 40060 42024 40069
rect 42340 40060 42392 40112
rect 42984 40128 43036 40180
rect 42524 39924 42576 39976
rect 43168 39992 43220 40044
rect 45284 40128 45336 40180
rect 47492 40128 47544 40180
rect 48320 40060 48372 40112
rect 44456 39992 44508 40044
rect 47032 39992 47084 40044
rect 49516 40060 49568 40112
rect 53380 40060 53432 40112
rect 53564 40060 53616 40112
rect 53932 40128 53984 40180
rect 54116 40128 54168 40180
rect 54668 40128 54720 40180
rect 57244 40128 57296 40180
rect 50252 39992 50304 40044
rect 52092 39992 52144 40044
rect 53656 39992 53708 40044
rect 54116 39992 54168 40044
rect 54484 39992 54536 40044
rect 55680 40060 55732 40112
rect 56600 39992 56652 40044
rect 57244 39992 57296 40044
rect 43536 39924 43588 39976
rect 48320 39924 48372 39976
rect 38108 39831 38160 39840
rect 38108 39797 38117 39831
rect 38117 39797 38151 39831
rect 38151 39797 38160 39831
rect 38108 39788 38160 39797
rect 46664 39856 46716 39908
rect 52920 39924 52972 39976
rect 54852 39967 54904 39976
rect 54852 39933 54861 39967
rect 54861 39933 54895 39967
rect 54895 39933 54904 39967
rect 54852 39924 54904 39933
rect 49608 39856 49660 39908
rect 50160 39856 50212 39908
rect 53196 39899 53248 39908
rect 53196 39865 53205 39899
rect 53205 39865 53239 39899
rect 53239 39865 53248 39899
rect 53196 39856 53248 39865
rect 53564 39856 53616 39908
rect 43904 39788 43956 39840
rect 47676 39788 47728 39840
rect 51724 39788 51776 39840
rect 53380 39788 53432 39840
rect 55588 39788 55640 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 29000 39627 29052 39636
rect 29000 39593 29009 39627
rect 29009 39593 29043 39627
rect 29043 39593 29052 39627
rect 29000 39584 29052 39593
rect 30656 39584 30708 39636
rect 31392 39584 31444 39636
rect 31852 39584 31904 39636
rect 32588 39627 32640 39636
rect 32588 39593 32597 39627
rect 32597 39593 32631 39627
rect 32631 39593 32640 39627
rect 32588 39584 32640 39593
rect 34060 39627 34112 39636
rect 34060 39593 34069 39627
rect 34069 39593 34103 39627
rect 34103 39593 34112 39627
rect 34060 39584 34112 39593
rect 36084 39627 36136 39636
rect 36084 39593 36093 39627
rect 36093 39593 36127 39627
rect 36127 39593 36136 39627
rect 36084 39584 36136 39593
rect 37004 39627 37056 39636
rect 37004 39593 37013 39627
rect 37013 39593 37047 39627
rect 37047 39593 37056 39627
rect 37004 39584 37056 39593
rect 30564 39516 30616 39568
rect 29184 39491 29236 39500
rect 29184 39457 29193 39491
rect 29193 39457 29227 39491
rect 29227 39457 29236 39491
rect 29184 39448 29236 39457
rect 33876 39491 33928 39500
rect 33876 39457 33885 39491
rect 33885 39457 33919 39491
rect 33919 39457 33928 39491
rect 33876 39448 33928 39457
rect 35256 39448 35308 39500
rect 37648 39516 37700 39568
rect 37740 39516 37792 39568
rect 38292 39516 38344 39568
rect 39948 39516 40000 39568
rect 40408 39516 40460 39568
rect 40684 39516 40736 39568
rect 29828 39423 29880 39432
rect 29828 39389 29837 39423
rect 29837 39389 29871 39423
rect 29871 39389 29880 39423
rect 29828 39380 29880 39389
rect 30656 39380 30708 39432
rect 33508 39380 33560 39432
rect 35440 39423 35492 39432
rect 35440 39389 35449 39423
rect 35449 39389 35483 39423
rect 35483 39389 35492 39423
rect 35440 39380 35492 39389
rect 35532 39423 35584 39432
rect 35532 39389 35542 39423
rect 35542 39389 35576 39423
rect 35576 39389 35584 39423
rect 37832 39448 37884 39500
rect 38108 39491 38160 39500
rect 38108 39457 38117 39491
rect 38117 39457 38151 39491
rect 38151 39457 38160 39491
rect 38108 39448 38160 39457
rect 38844 39491 38896 39500
rect 38844 39457 38853 39491
rect 38853 39457 38887 39491
rect 38887 39457 38896 39491
rect 38844 39448 38896 39457
rect 40960 39448 41012 39500
rect 35532 39380 35584 39389
rect 35992 39380 36044 39432
rect 36912 39380 36964 39432
rect 30380 39312 30432 39364
rect 30564 39312 30616 39364
rect 31392 39355 31444 39364
rect 31392 39321 31401 39355
rect 31401 39321 31435 39355
rect 31435 39321 31444 39355
rect 31392 39312 31444 39321
rect 32312 39355 32364 39364
rect 32312 39321 32321 39355
rect 32321 39321 32355 39355
rect 32355 39321 32364 39355
rect 32312 39312 32364 39321
rect 34796 39312 34848 39364
rect 39580 39380 39632 39432
rect 39856 39380 39908 39432
rect 42156 39516 42208 39568
rect 34428 39244 34480 39296
rect 39672 39312 39724 39364
rect 42064 39423 42116 39432
rect 42524 39448 42576 39500
rect 42064 39389 42109 39423
rect 42109 39389 42116 39423
rect 42064 39380 42116 39389
rect 42708 39423 42760 39432
rect 42708 39389 42717 39423
rect 42717 39389 42751 39423
rect 42751 39389 42760 39423
rect 42708 39380 42760 39389
rect 42800 39423 42852 39432
rect 42800 39389 42837 39423
rect 42837 39389 42852 39423
rect 42800 39380 42852 39389
rect 43168 39423 43220 39432
rect 43168 39389 43182 39423
rect 43182 39389 43216 39423
rect 43216 39389 43220 39423
rect 44272 39423 44324 39432
rect 43168 39380 43220 39389
rect 44272 39389 44281 39423
rect 44281 39389 44315 39423
rect 44315 39389 44324 39423
rect 44272 39380 44324 39389
rect 46940 39423 46992 39432
rect 41880 39355 41932 39364
rect 36912 39244 36964 39296
rect 41420 39244 41472 39296
rect 41880 39321 41889 39355
rect 41889 39321 41923 39355
rect 41923 39321 41932 39355
rect 41880 39312 41932 39321
rect 42984 39355 43036 39364
rect 42984 39321 42993 39355
rect 42993 39321 43027 39355
rect 43027 39321 43036 39355
rect 42984 39312 43036 39321
rect 45560 39312 45612 39364
rect 42432 39244 42484 39296
rect 45468 39244 45520 39296
rect 46940 39389 46949 39423
rect 46949 39389 46983 39423
rect 46983 39389 46992 39423
rect 46940 39380 46992 39389
rect 47032 39423 47084 39432
rect 47032 39389 47041 39423
rect 47041 39389 47075 39423
rect 47075 39389 47084 39423
rect 49792 39516 49844 39568
rect 52092 39516 52144 39568
rect 47032 39380 47084 39389
rect 49700 39448 49752 39500
rect 51724 39448 51776 39500
rect 48504 39423 48556 39432
rect 48504 39389 48518 39423
rect 48518 39389 48552 39423
rect 48552 39389 48556 39423
rect 48504 39380 48556 39389
rect 48872 39380 48924 39432
rect 47216 39355 47268 39364
rect 47216 39321 47225 39355
rect 47225 39321 47259 39355
rect 47259 39321 47268 39355
rect 47216 39312 47268 39321
rect 48320 39355 48372 39364
rect 48320 39321 48329 39355
rect 48329 39321 48363 39355
rect 48363 39321 48372 39355
rect 48320 39312 48372 39321
rect 48412 39355 48464 39364
rect 48412 39321 48421 39355
rect 48421 39321 48455 39355
rect 48455 39321 48464 39355
rect 48412 39312 48464 39321
rect 48136 39244 48188 39296
rect 50988 39312 51040 39364
rect 48688 39244 48740 39296
rect 49332 39244 49384 39296
rect 51632 39355 51684 39364
rect 51632 39321 51641 39355
rect 51641 39321 51675 39355
rect 51675 39321 51684 39355
rect 51632 39312 51684 39321
rect 51816 39380 51868 39432
rect 51724 39287 51776 39296
rect 51724 39253 51739 39287
rect 51739 39253 51773 39287
rect 51773 39253 51776 39287
rect 51724 39244 51776 39253
rect 51908 39244 51960 39296
rect 53380 39491 53432 39500
rect 53380 39457 53389 39491
rect 53389 39457 53423 39491
rect 53423 39457 53432 39491
rect 53380 39448 53432 39457
rect 53748 39448 53800 39500
rect 55956 39448 56008 39500
rect 54116 39423 54168 39432
rect 54116 39389 54126 39423
rect 54126 39389 54160 39423
rect 54160 39389 54168 39423
rect 54116 39380 54168 39389
rect 54300 39423 54352 39432
rect 54300 39389 54309 39423
rect 54309 39389 54343 39423
rect 54343 39389 54352 39423
rect 54300 39380 54352 39389
rect 54760 39380 54812 39432
rect 55772 39423 55824 39432
rect 55772 39389 55781 39423
rect 55781 39389 55815 39423
rect 55815 39389 55824 39423
rect 55772 39380 55824 39389
rect 56876 39380 56928 39432
rect 57244 39423 57296 39432
rect 57244 39389 57253 39423
rect 57253 39389 57287 39423
rect 57287 39389 57296 39423
rect 57244 39380 57296 39389
rect 55588 39312 55640 39364
rect 53472 39244 53524 39296
rect 54116 39244 54168 39296
rect 56048 39244 56100 39296
rect 56508 39244 56560 39296
rect 58440 39244 58492 39296
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 35594 39142 35646 39194
rect 35658 39142 35710 39194
rect 35722 39142 35774 39194
rect 35786 39142 35838 39194
rect 35850 39142 35902 39194
rect 30564 39083 30616 39092
rect 30564 39049 30573 39083
rect 30573 39049 30607 39083
rect 30607 39049 30616 39083
rect 30564 39040 30616 39049
rect 31668 39040 31720 39092
rect 32496 39040 32548 39092
rect 34428 39083 34480 39092
rect 29736 38947 29788 38956
rect 29736 38913 29745 38947
rect 29745 38913 29779 38947
rect 29779 38913 29788 38947
rect 29736 38904 29788 38913
rect 30840 38904 30892 38956
rect 32772 38972 32824 39024
rect 34428 39049 34437 39083
rect 34437 39049 34471 39083
rect 34471 39049 34480 39083
rect 34428 39040 34480 39049
rect 35440 39040 35492 39092
rect 44272 39040 44324 39092
rect 47032 39040 47084 39092
rect 47584 39040 47636 39092
rect 36544 39015 36596 39024
rect 29184 38836 29236 38888
rect 32312 38904 32364 38956
rect 32680 38904 32732 38956
rect 33600 38904 33652 38956
rect 34612 38904 34664 38956
rect 35256 38947 35308 38956
rect 35256 38913 35265 38947
rect 35265 38913 35299 38947
rect 35299 38913 35308 38947
rect 35256 38904 35308 38913
rect 36544 38981 36553 39015
rect 36553 38981 36587 39015
rect 36587 38981 36596 39015
rect 36544 38972 36596 38981
rect 41420 38972 41472 39024
rect 42432 38972 42484 39024
rect 33876 38836 33928 38888
rect 34704 38836 34756 38888
rect 35348 38879 35400 38888
rect 35348 38845 35357 38879
rect 35357 38845 35391 38879
rect 35391 38845 35400 38879
rect 35348 38836 35400 38845
rect 35440 38836 35492 38888
rect 33048 38768 33100 38820
rect 36820 38947 36872 38956
rect 36820 38913 36828 38947
rect 36828 38913 36862 38947
rect 36862 38913 36872 38947
rect 36820 38904 36872 38913
rect 36912 38947 36964 38956
rect 36912 38913 36921 38947
rect 36921 38913 36955 38947
rect 36955 38913 36964 38947
rect 36912 38904 36964 38913
rect 38108 38904 38160 38956
rect 38660 38904 38712 38956
rect 40040 38904 40092 38956
rect 42892 38947 42944 38956
rect 39856 38879 39908 38888
rect 39856 38845 39865 38879
rect 39865 38845 39899 38879
rect 39899 38845 39908 38879
rect 39856 38836 39908 38845
rect 41052 38879 41104 38888
rect 41052 38845 41061 38879
rect 41061 38845 41095 38879
rect 41095 38845 41104 38879
rect 41052 38836 41104 38845
rect 37740 38768 37792 38820
rect 41972 38836 42024 38888
rect 42892 38913 42901 38947
rect 42901 38913 42935 38947
rect 42935 38913 42944 38947
rect 42892 38904 42944 38913
rect 42800 38836 42852 38888
rect 43168 38904 43220 38956
rect 44180 38947 44232 38956
rect 44180 38913 44189 38947
rect 44189 38913 44223 38947
rect 44223 38913 44232 38947
rect 44180 38904 44232 38913
rect 45008 38947 45060 38956
rect 45008 38913 45017 38947
rect 45017 38913 45051 38947
rect 45051 38913 45060 38947
rect 45008 38904 45060 38913
rect 45192 38947 45244 38956
rect 45192 38913 45201 38947
rect 45201 38913 45235 38947
rect 45235 38913 45244 38947
rect 45192 38904 45244 38913
rect 48412 39040 48464 39092
rect 48136 38972 48188 39024
rect 48320 38947 48372 38956
rect 48320 38913 48329 38947
rect 48329 38913 48363 38947
rect 48363 38913 48372 38947
rect 48320 38904 48372 38913
rect 48872 39040 48924 39092
rect 55772 39040 55824 39092
rect 56876 39083 56928 39092
rect 56876 39049 56885 39083
rect 56885 39049 56919 39083
rect 56919 39049 56928 39083
rect 56876 39040 56928 39049
rect 47216 38836 47268 38888
rect 47768 38836 47820 38888
rect 47860 38836 47912 38888
rect 30380 38700 30432 38752
rect 32220 38700 32272 38752
rect 37280 38700 37332 38752
rect 37556 38743 37608 38752
rect 37556 38709 37565 38743
rect 37565 38709 37599 38743
rect 37599 38709 37608 38743
rect 37556 38700 37608 38709
rect 42064 38700 42116 38752
rect 42708 38700 42760 38752
rect 45744 38768 45796 38820
rect 47124 38768 47176 38820
rect 43812 38700 43864 38752
rect 45652 38743 45704 38752
rect 45652 38709 45661 38743
rect 45661 38709 45695 38743
rect 45695 38709 45704 38743
rect 45652 38700 45704 38709
rect 47860 38743 47912 38752
rect 47860 38709 47869 38743
rect 47869 38709 47903 38743
rect 47903 38709 47912 38743
rect 47860 38700 47912 38709
rect 51632 38972 51684 39024
rect 51724 38972 51776 39024
rect 49056 38904 49108 38956
rect 50712 38904 50764 38956
rect 51080 38947 51132 38956
rect 51080 38913 51089 38947
rect 51089 38913 51123 38947
rect 51123 38913 51132 38947
rect 51080 38904 51132 38913
rect 52000 38904 52052 38956
rect 52828 38904 52880 38956
rect 53472 38947 53524 38956
rect 51172 38879 51224 38888
rect 51172 38845 51181 38879
rect 51181 38845 51215 38879
rect 51215 38845 51224 38879
rect 51172 38836 51224 38845
rect 50804 38768 50856 38820
rect 51816 38768 51868 38820
rect 49332 38700 49384 38752
rect 50344 38700 50396 38752
rect 52000 38768 52052 38820
rect 52276 38768 52328 38820
rect 53472 38913 53480 38947
rect 53480 38913 53514 38947
rect 53514 38913 53524 38947
rect 53472 38904 53524 38913
rect 54116 38972 54168 39024
rect 54208 38947 54260 38956
rect 54208 38913 54217 38947
rect 54217 38913 54251 38947
rect 54251 38913 54260 38947
rect 54208 38904 54260 38913
rect 54392 38972 54444 39024
rect 53840 38836 53892 38888
rect 54024 38836 54076 38888
rect 54668 38947 54720 38956
rect 54668 38913 54682 38947
rect 54682 38913 54716 38947
rect 54716 38913 54720 38947
rect 56508 38947 56560 38956
rect 54668 38904 54720 38913
rect 56508 38913 56517 38947
rect 56517 38913 56551 38947
rect 56551 38913 56560 38947
rect 56508 38904 56560 38913
rect 56048 38836 56100 38888
rect 52736 38700 52788 38752
rect 53012 38700 53064 38752
rect 55220 38700 55272 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 30656 38496 30708 38548
rect 33876 38539 33928 38548
rect 31852 38428 31904 38480
rect 30104 38292 30156 38344
rect 30380 38292 30432 38344
rect 29736 38224 29788 38276
rect 30748 38156 30800 38208
rect 31208 38292 31260 38344
rect 32220 38335 32272 38344
rect 32220 38301 32229 38335
rect 32229 38301 32263 38335
rect 32263 38301 32272 38335
rect 32220 38292 32272 38301
rect 31576 38224 31628 38276
rect 31668 38224 31720 38276
rect 33876 38505 33885 38539
rect 33885 38505 33919 38539
rect 33919 38505 33928 38539
rect 33876 38496 33928 38505
rect 35348 38539 35400 38548
rect 35348 38505 35357 38539
rect 35357 38505 35391 38539
rect 35391 38505 35400 38539
rect 35348 38496 35400 38505
rect 35440 38496 35492 38548
rect 41052 38539 41104 38548
rect 41052 38505 41061 38539
rect 41061 38505 41095 38539
rect 41095 38505 41104 38539
rect 41052 38496 41104 38505
rect 47216 38539 47268 38548
rect 47216 38505 47225 38539
rect 47225 38505 47259 38539
rect 47259 38505 47268 38539
rect 47216 38496 47268 38505
rect 48320 38496 48372 38548
rect 51080 38496 51132 38548
rect 51908 38496 51960 38548
rect 52920 38496 52972 38548
rect 53472 38496 53524 38548
rect 54208 38496 54260 38548
rect 55312 38496 55364 38548
rect 55588 38496 55640 38548
rect 32496 38335 32548 38344
rect 32496 38301 32505 38335
rect 32505 38301 32539 38335
rect 32539 38301 32548 38335
rect 32496 38292 32548 38301
rect 32680 38335 32732 38344
rect 32680 38301 32694 38335
rect 32694 38301 32728 38335
rect 32728 38301 32732 38335
rect 34612 38428 34664 38480
rect 33416 38403 33468 38412
rect 33416 38369 33425 38403
rect 33425 38369 33459 38403
rect 33459 38369 33468 38403
rect 33416 38360 33468 38369
rect 33692 38360 33744 38412
rect 36728 38428 36780 38480
rect 32680 38292 32732 38301
rect 34520 38292 34572 38344
rect 35072 38335 35124 38344
rect 35072 38301 35081 38335
rect 35081 38301 35115 38335
rect 35115 38301 35124 38335
rect 35072 38292 35124 38301
rect 34980 38224 35032 38276
rect 36360 38292 36412 38344
rect 36636 38335 36688 38344
rect 36636 38301 36645 38335
rect 36645 38301 36679 38335
rect 36679 38301 36688 38335
rect 36636 38292 36688 38301
rect 36820 38335 36872 38344
rect 36820 38301 36829 38335
rect 36829 38301 36863 38335
rect 36863 38301 36872 38335
rect 36820 38292 36872 38301
rect 37280 38292 37332 38344
rect 40040 38428 40092 38480
rect 44180 38428 44232 38480
rect 38660 38360 38712 38412
rect 37924 38335 37976 38344
rect 37924 38301 37933 38335
rect 37933 38301 37967 38335
rect 37967 38301 37976 38335
rect 37924 38292 37976 38301
rect 38108 38292 38160 38344
rect 40132 38360 40184 38412
rect 39488 38292 39540 38344
rect 39764 38292 39816 38344
rect 41880 38360 41932 38412
rect 42524 38360 42576 38412
rect 45744 38403 45796 38412
rect 45744 38369 45753 38403
rect 45753 38369 45787 38403
rect 45787 38369 45796 38403
rect 45744 38360 45796 38369
rect 47216 38360 47268 38412
rect 49056 38360 49108 38412
rect 49240 38403 49292 38412
rect 49240 38369 49249 38403
rect 49249 38369 49283 38403
rect 49283 38369 49292 38403
rect 49240 38360 49292 38369
rect 51172 38428 51224 38480
rect 53840 38428 53892 38480
rect 54852 38428 54904 38480
rect 40684 38335 40736 38344
rect 40684 38301 40693 38335
rect 40693 38301 40727 38335
rect 40727 38301 40736 38335
rect 40684 38292 40736 38301
rect 40960 38292 41012 38344
rect 43536 38335 43588 38344
rect 43536 38301 43545 38335
rect 43545 38301 43579 38335
rect 43579 38301 43588 38335
rect 43536 38292 43588 38301
rect 45560 38335 45612 38344
rect 45560 38301 45569 38335
rect 45569 38301 45603 38335
rect 45603 38301 45612 38335
rect 45560 38292 45612 38301
rect 46940 38292 46992 38344
rect 49424 38292 49476 38344
rect 50344 38335 50396 38344
rect 50344 38301 50353 38335
rect 50353 38301 50387 38335
rect 50387 38301 50396 38335
rect 50344 38292 50396 38301
rect 50436 38335 50488 38344
rect 50436 38301 50446 38335
rect 50446 38301 50480 38335
rect 50480 38301 50488 38335
rect 50436 38292 50488 38301
rect 50804 38335 50856 38344
rect 50804 38301 50818 38335
rect 50818 38301 50852 38335
rect 50852 38301 50856 38335
rect 53012 38360 53064 38412
rect 53564 38360 53616 38412
rect 54208 38360 54260 38412
rect 55220 38360 55272 38412
rect 50804 38292 50856 38301
rect 53196 38292 53248 38344
rect 31852 38156 31904 38208
rect 35072 38156 35124 38208
rect 40224 38224 40276 38276
rect 36728 38199 36780 38208
rect 36728 38165 36737 38199
rect 36737 38165 36771 38199
rect 36771 38165 36780 38199
rect 36728 38156 36780 38165
rect 37832 38156 37884 38208
rect 39580 38156 39632 38208
rect 40408 38156 40460 38208
rect 42340 38224 42392 38276
rect 42432 38224 42484 38276
rect 42800 38224 42852 38276
rect 47768 38224 47820 38276
rect 42156 38156 42208 38208
rect 45652 38156 45704 38208
rect 47676 38156 47728 38208
rect 48688 38199 48740 38208
rect 48688 38165 48697 38199
rect 48697 38165 48731 38199
rect 48731 38165 48740 38199
rect 48688 38156 48740 38165
rect 50712 38267 50764 38276
rect 50712 38233 50721 38267
rect 50721 38233 50755 38267
rect 50755 38233 50764 38267
rect 50712 38224 50764 38233
rect 50896 38224 50948 38276
rect 52368 38224 52420 38276
rect 54024 38292 54076 38344
rect 55680 38335 55732 38344
rect 55680 38301 55689 38335
rect 55689 38301 55723 38335
rect 55723 38301 55732 38335
rect 55680 38292 55732 38301
rect 52000 38156 52052 38208
rect 54484 38156 54536 38208
rect 56048 38199 56100 38208
rect 56048 38165 56057 38199
rect 56057 38165 56091 38199
rect 56091 38165 56100 38199
rect 56048 38156 56100 38165
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 35594 38054 35646 38106
rect 35658 38054 35710 38106
rect 35722 38054 35774 38106
rect 35786 38054 35838 38106
rect 35850 38054 35902 38106
rect 29276 37995 29328 38004
rect 29276 37961 29285 37995
rect 29285 37961 29319 37995
rect 29319 37961 29328 37995
rect 29276 37952 29328 37961
rect 31484 37952 31536 38004
rect 33048 37952 33100 38004
rect 29184 37859 29236 37868
rect 29184 37825 29193 37859
rect 29193 37825 29227 37859
rect 29227 37825 29236 37859
rect 29184 37816 29236 37825
rect 30564 37884 30616 37936
rect 31944 37884 31996 37936
rect 32496 37927 32548 37936
rect 32496 37893 32505 37927
rect 32505 37893 32539 37927
rect 32539 37893 32548 37927
rect 34796 37952 34848 38004
rect 32496 37884 32548 37893
rect 33508 37884 33560 37936
rect 33692 37884 33744 37936
rect 30380 37816 30432 37868
rect 30932 37859 30984 37868
rect 30196 37791 30248 37800
rect 30196 37757 30205 37791
rect 30205 37757 30239 37791
rect 30239 37757 30248 37791
rect 30196 37748 30248 37757
rect 30932 37825 30941 37859
rect 30941 37825 30975 37859
rect 30975 37825 30984 37859
rect 30932 37816 30984 37825
rect 31208 37816 31260 37868
rect 31576 37816 31628 37868
rect 35532 37884 35584 37936
rect 35992 37927 36044 37936
rect 30840 37748 30892 37800
rect 29276 37612 29328 37664
rect 33784 37612 33836 37664
rect 34980 37816 35032 37868
rect 35440 37816 35492 37868
rect 35992 37893 36001 37927
rect 36001 37893 36035 37927
rect 36035 37893 36044 37927
rect 35992 37884 36044 37893
rect 38936 37952 38988 38004
rect 39488 37952 39540 38004
rect 39764 37995 39816 38004
rect 39764 37961 39773 37995
rect 39773 37961 39807 37995
rect 39807 37961 39816 37995
rect 39764 37952 39816 37961
rect 40776 37952 40828 38004
rect 41696 37952 41748 38004
rect 41880 37952 41932 38004
rect 42248 37952 42300 38004
rect 36360 37816 36412 37868
rect 36636 37859 36688 37868
rect 36636 37825 36645 37859
rect 36645 37825 36679 37859
rect 36679 37825 36688 37859
rect 36636 37816 36688 37825
rect 37832 37816 37884 37868
rect 39488 37859 39540 37868
rect 39488 37825 39497 37859
rect 39497 37825 39531 37859
rect 39531 37825 39540 37859
rect 39488 37816 39540 37825
rect 39672 37816 39724 37868
rect 40224 37884 40276 37936
rect 42892 37927 42944 37936
rect 40408 37816 40460 37868
rect 42892 37893 42901 37927
rect 42901 37893 42935 37927
rect 42935 37893 42944 37927
rect 42892 37884 42944 37893
rect 51908 37952 51960 38004
rect 52368 37952 52420 38004
rect 54116 37952 54168 38004
rect 54852 37952 54904 38004
rect 43812 37927 43864 37936
rect 43812 37893 43821 37927
rect 43821 37893 43855 37927
rect 43855 37893 43864 37927
rect 43812 37884 43864 37893
rect 45284 37884 45336 37936
rect 42616 37859 42668 37868
rect 42616 37825 42625 37859
rect 42625 37825 42659 37859
rect 42659 37825 42668 37859
rect 42616 37816 42668 37825
rect 42708 37859 42760 37868
rect 42708 37825 42718 37859
rect 42718 37825 42752 37859
rect 42752 37825 42760 37859
rect 42708 37816 42760 37825
rect 43076 37859 43128 37868
rect 43076 37825 43090 37859
rect 43090 37825 43124 37859
rect 43124 37825 43128 37859
rect 43076 37816 43128 37825
rect 42064 37748 42116 37800
rect 42524 37748 42576 37800
rect 43720 37748 43772 37800
rect 39948 37680 40000 37732
rect 41696 37680 41748 37732
rect 48320 37884 48372 37936
rect 48688 37884 48740 37936
rect 49332 37884 49384 37936
rect 56140 37884 56192 37936
rect 46112 37816 46164 37868
rect 46940 37859 46992 37868
rect 46020 37748 46072 37800
rect 46940 37825 46949 37859
rect 46949 37825 46983 37859
rect 46983 37825 46992 37859
rect 46940 37816 46992 37825
rect 47768 37816 47820 37868
rect 48228 37859 48280 37868
rect 48228 37825 48238 37859
rect 48238 37825 48272 37859
rect 48272 37825 48280 37859
rect 48228 37816 48280 37825
rect 48412 37859 48464 37868
rect 48412 37825 48421 37859
rect 48421 37825 48455 37859
rect 48455 37825 48464 37859
rect 48412 37816 48464 37825
rect 48596 37859 48648 37868
rect 48596 37825 48610 37859
rect 48610 37825 48644 37859
rect 48644 37825 48648 37859
rect 48596 37816 48648 37825
rect 53196 37859 53248 37868
rect 53196 37825 53205 37859
rect 53205 37825 53239 37859
rect 53239 37825 53248 37859
rect 53196 37816 53248 37825
rect 55956 37859 56008 37868
rect 55956 37825 55965 37859
rect 55965 37825 55999 37859
rect 55999 37825 56008 37859
rect 55956 37816 56008 37825
rect 56324 37816 56376 37868
rect 50804 37791 50856 37800
rect 35348 37612 35400 37664
rect 37556 37612 37608 37664
rect 39488 37612 39540 37664
rect 40408 37612 40460 37664
rect 40776 37612 40828 37664
rect 41972 37612 42024 37664
rect 43352 37612 43404 37664
rect 46480 37655 46532 37664
rect 46480 37621 46489 37655
rect 46489 37621 46523 37655
rect 46523 37621 46532 37655
rect 46480 37612 46532 37621
rect 50804 37757 50813 37791
rect 50813 37757 50847 37791
rect 50847 37757 50856 37791
rect 50804 37748 50856 37757
rect 54484 37748 54536 37800
rect 55864 37791 55916 37800
rect 55864 37757 55873 37791
rect 55873 37757 55907 37791
rect 55907 37757 55916 37791
rect 55864 37748 55916 37757
rect 56048 37748 56100 37800
rect 57704 37680 57756 37732
rect 49792 37655 49844 37664
rect 49792 37621 49801 37655
rect 49801 37621 49835 37655
rect 49835 37621 49844 37655
rect 49792 37612 49844 37621
rect 50436 37612 50488 37664
rect 50896 37612 50948 37664
rect 57244 37655 57296 37664
rect 57244 37621 57253 37655
rect 57253 37621 57287 37655
rect 57287 37621 57296 37655
rect 57244 37612 57296 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 30656 37408 30708 37460
rect 32312 37451 32364 37460
rect 32312 37417 32321 37451
rect 32321 37417 32355 37451
rect 32355 37417 32364 37451
rect 32312 37408 32364 37417
rect 32680 37408 32732 37460
rect 32772 37408 32824 37460
rect 37464 37408 37516 37460
rect 37648 37408 37700 37460
rect 38108 37408 38160 37460
rect 28172 37247 28224 37256
rect 28172 37213 28181 37247
rect 28181 37213 28215 37247
rect 28215 37213 28224 37247
rect 28172 37204 28224 37213
rect 34060 37340 34112 37392
rect 35624 37383 35676 37392
rect 35624 37349 35633 37383
rect 35633 37349 35667 37383
rect 35667 37349 35676 37383
rect 35624 37340 35676 37349
rect 28816 37272 28868 37324
rect 29368 37272 29420 37324
rect 30748 37315 30800 37324
rect 30748 37281 30757 37315
rect 30757 37281 30791 37315
rect 30791 37281 30800 37315
rect 30748 37272 30800 37281
rect 30932 37315 30984 37324
rect 30932 37281 30941 37315
rect 30941 37281 30975 37315
rect 30975 37281 30984 37315
rect 30932 37272 30984 37281
rect 32680 37272 32732 37324
rect 33876 37272 33928 37324
rect 36636 37340 36688 37392
rect 39672 37340 39724 37392
rect 42616 37408 42668 37460
rect 43720 37451 43772 37460
rect 43720 37417 43729 37451
rect 43729 37417 43763 37451
rect 43763 37417 43772 37451
rect 43720 37408 43772 37417
rect 46940 37408 46992 37460
rect 52460 37408 52512 37460
rect 53472 37451 53524 37460
rect 53472 37417 53481 37451
rect 53481 37417 53515 37451
rect 53515 37417 53524 37451
rect 53472 37408 53524 37417
rect 56324 37451 56376 37460
rect 56324 37417 56333 37451
rect 56333 37417 56367 37451
rect 56367 37417 56376 37451
rect 56324 37408 56376 37417
rect 40684 37340 40736 37392
rect 30564 37247 30616 37256
rect 30564 37213 30573 37247
rect 30573 37213 30607 37247
rect 30607 37213 30616 37247
rect 30564 37204 30616 37213
rect 28264 37111 28316 37120
rect 28264 37077 28273 37111
rect 28273 37077 28307 37111
rect 28307 37077 28316 37111
rect 28264 37068 28316 37077
rect 29276 37136 29328 37188
rect 30196 37136 30248 37188
rect 32956 37136 33008 37188
rect 28908 37068 28960 37120
rect 29092 37068 29144 37120
rect 33140 37136 33192 37188
rect 33508 37204 33560 37256
rect 33692 37204 33744 37256
rect 34612 37204 34664 37256
rect 33784 37179 33836 37188
rect 33784 37145 33793 37179
rect 33793 37145 33827 37179
rect 33827 37145 33836 37179
rect 33784 37136 33836 37145
rect 33876 37136 33928 37188
rect 35992 37204 36044 37256
rect 36728 37272 36780 37324
rect 38384 37272 38436 37324
rect 36360 37247 36412 37256
rect 36360 37213 36369 37247
rect 36369 37213 36403 37247
rect 36403 37213 36412 37247
rect 36360 37204 36412 37213
rect 36636 37247 36688 37256
rect 36636 37213 36645 37247
rect 36645 37213 36679 37247
rect 36679 37213 36688 37247
rect 36636 37204 36688 37213
rect 37740 37204 37792 37256
rect 39028 37315 39080 37324
rect 39028 37281 39037 37315
rect 39037 37281 39071 37315
rect 39071 37281 39080 37315
rect 39028 37272 39080 37281
rect 39580 37272 39632 37324
rect 43352 37315 43404 37324
rect 40040 37247 40092 37256
rect 40040 37213 40049 37247
rect 40049 37213 40083 37247
rect 40083 37213 40092 37247
rect 40040 37204 40092 37213
rect 34428 37068 34480 37120
rect 39212 37136 39264 37188
rect 39948 37136 40000 37188
rect 40592 37204 40644 37256
rect 41512 37247 41564 37256
rect 41512 37213 41521 37247
rect 41521 37213 41555 37247
rect 41555 37213 41564 37247
rect 41512 37204 41564 37213
rect 41788 37247 41840 37256
rect 41788 37213 41797 37247
rect 41797 37213 41831 37247
rect 41831 37213 41840 37247
rect 41788 37204 41840 37213
rect 42248 37247 42300 37256
rect 42248 37213 42257 37247
rect 42257 37213 42291 37247
rect 42291 37213 42300 37247
rect 43352 37281 43361 37315
rect 43361 37281 43395 37315
rect 43395 37281 43404 37315
rect 43352 37272 43404 37281
rect 42248 37204 42300 37213
rect 43444 37247 43496 37256
rect 43444 37213 43453 37247
rect 43453 37213 43487 37247
rect 43487 37213 43496 37247
rect 43444 37204 43496 37213
rect 46020 37247 46072 37256
rect 46020 37213 46029 37247
rect 46029 37213 46063 37247
rect 46063 37213 46072 37247
rect 46020 37204 46072 37213
rect 46112 37204 46164 37256
rect 46572 37204 46624 37256
rect 46940 37204 46992 37256
rect 49332 37340 49384 37392
rect 52000 37340 52052 37392
rect 52920 37340 52972 37392
rect 48596 37272 48648 37324
rect 50252 37272 50304 37324
rect 53288 37272 53340 37324
rect 42708 37136 42760 37188
rect 35624 37068 35676 37120
rect 37464 37068 37516 37120
rect 37832 37111 37884 37120
rect 37832 37077 37841 37111
rect 37841 37077 37875 37111
rect 37875 37077 37884 37111
rect 37832 37068 37884 37077
rect 42524 37068 42576 37120
rect 45008 37068 45060 37120
rect 45100 37068 45152 37120
rect 45468 37068 45520 37120
rect 48320 37247 48372 37256
rect 48320 37213 48330 37247
rect 48330 37213 48364 37247
rect 48364 37213 48372 37247
rect 48320 37204 48372 37213
rect 49332 37247 49384 37256
rect 49332 37213 49341 37247
rect 49341 37213 49375 37247
rect 49375 37213 49384 37247
rect 49332 37204 49384 37213
rect 47768 37179 47820 37188
rect 47768 37145 47777 37179
rect 47777 37145 47811 37179
rect 47811 37145 47820 37179
rect 47768 37136 47820 37145
rect 48412 37136 48464 37188
rect 49700 37204 49752 37256
rect 50804 37204 50856 37256
rect 50988 37204 51040 37256
rect 54116 37340 54168 37392
rect 54484 37340 54536 37392
rect 53564 37272 53616 37324
rect 47860 37068 47912 37120
rect 50344 37136 50396 37188
rect 52460 37136 52512 37188
rect 48688 37068 48740 37120
rect 49148 37068 49200 37120
rect 52000 37068 52052 37120
rect 53196 37068 53248 37120
rect 54208 37247 54260 37256
rect 54208 37213 54218 37247
rect 54218 37213 54252 37247
rect 54252 37213 54260 37247
rect 55864 37272 55916 37324
rect 54208 37204 54260 37213
rect 54576 37247 54628 37256
rect 54576 37213 54590 37247
rect 54590 37213 54624 37247
rect 54624 37213 54628 37247
rect 54576 37204 54628 37213
rect 55772 37204 55824 37256
rect 54392 37179 54444 37188
rect 54392 37145 54401 37179
rect 54401 37145 54435 37179
rect 54435 37145 54444 37179
rect 54392 37136 54444 37145
rect 54852 37068 54904 37120
rect 57980 37111 58032 37120
rect 57980 37077 57989 37111
rect 57989 37077 58023 37111
rect 58023 37077 58032 37111
rect 57980 37068 58032 37077
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 28264 36864 28316 36916
rect 29736 36864 29788 36916
rect 30012 36907 30064 36916
rect 30012 36873 30021 36907
rect 30021 36873 30055 36907
rect 30055 36873 30064 36907
rect 30012 36864 30064 36873
rect 33784 36864 33836 36916
rect 35808 36864 35860 36916
rect 36636 36864 36688 36916
rect 39028 36864 39080 36916
rect 39212 36864 39264 36916
rect 43536 36864 43588 36916
rect 30196 36796 30248 36848
rect 28172 36728 28224 36780
rect 28908 36771 28960 36780
rect 28908 36737 28917 36771
rect 28917 36737 28951 36771
rect 28951 36737 28960 36771
rect 28908 36728 28960 36737
rect 29092 36728 29144 36780
rect 29920 36771 29972 36780
rect 29920 36737 29929 36771
rect 29929 36737 29963 36771
rect 29963 36737 29972 36771
rect 29920 36728 29972 36737
rect 29368 36660 29420 36712
rect 30564 36728 30616 36780
rect 30932 36728 30984 36780
rect 31392 36796 31444 36848
rect 32864 36796 32916 36848
rect 32956 36796 33008 36848
rect 32680 36771 32732 36780
rect 32680 36737 32689 36771
rect 32689 36737 32723 36771
rect 32723 36737 32732 36771
rect 32680 36728 32732 36737
rect 32772 36728 32824 36780
rect 34428 36771 34480 36780
rect 34428 36737 34437 36771
rect 34437 36737 34471 36771
rect 34471 36737 34480 36771
rect 34428 36728 34480 36737
rect 34612 36728 34664 36780
rect 30380 36660 30432 36712
rect 30656 36703 30708 36712
rect 30656 36669 30665 36703
rect 30665 36669 30699 36703
rect 30699 36669 30708 36703
rect 30656 36660 30708 36669
rect 34244 36703 34296 36712
rect 34244 36669 34253 36703
rect 34253 36669 34287 36703
rect 34287 36669 34296 36703
rect 34244 36660 34296 36669
rect 29184 36635 29236 36644
rect 29184 36601 29193 36635
rect 29193 36601 29227 36635
rect 29227 36601 29236 36635
rect 29184 36592 29236 36601
rect 29276 36592 29328 36644
rect 33140 36524 33192 36576
rect 33968 36524 34020 36576
rect 37832 36796 37884 36848
rect 35992 36728 36044 36780
rect 35808 36660 35860 36712
rect 36176 36592 36228 36644
rect 37188 36728 37240 36780
rect 38108 36771 38160 36780
rect 38108 36737 38117 36771
rect 38117 36737 38151 36771
rect 38151 36737 38160 36771
rect 38108 36728 38160 36737
rect 38936 36771 38988 36780
rect 38936 36737 38945 36771
rect 38945 36737 38979 36771
rect 38979 36737 38988 36771
rect 38936 36728 38988 36737
rect 40040 36796 40092 36848
rect 38016 36703 38068 36712
rect 38016 36669 38025 36703
rect 38025 36669 38059 36703
rect 38059 36669 38068 36703
rect 38016 36660 38068 36669
rect 39212 36728 39264 36780
rect 39948 36728 40000 36780
rect 40224 36771 40276 36780
rect 40224 36737 40233 36771
rect 40233 36737 40267 36771
rect 40267 36737 40276 36771
rect 40224 36728 40276 36737
rect 41420 36771 41472 36780
rect 41420 36737 41429 36771
rect 41429 36737 41463 36771
rect 41463 36737 41472 36771
rect 41420 36728 41472 36737
rect 44088 36796 44140 36848
rect 42892 36771 42944 36780
rect 42892 36737 42901 36771
rect 42901 36737 42935 36771
rect 42935 36737 42944 36771
rect 42892 36728 42944 36737
rect 44272 36728 44324 36780
rect 45192 36728 45244 36780
rect 45468 36771 45520 36780
rect 45468 36737 45477 36771
rect 45477 36737 45511 36771
rect 45511 36737 45520 36771
rect 45468 36728 45520 36737
rect 47768 36796 47820 36848
rect 48596 36864 48648 36916
rect 50068 36864 50120 36916
rect 50712 36864 50764 36916
rect 49976 36796 50028 36848
rect 50344 36839 50396 36848
rect 50344 36805 50353 36839
rect 50353 36805 50387 36839
rect 50387 36805 50396 36839
rect 50344 36796 50396 36805
rect 52368 36864 52420 36916
rect 52920 36864 52972 36916
rect 52000 36796 52052 36848
rect 46020 36728 46072 36780
rect 46296 36728 46348 36780
rect 46572 36728 46624 36780
rect 49240 36771 49292 36780
rect 49240 36737 49249 36771
rect 49249 36737 49283 36771
rect 49283 36737 49292 36771
rect 49240 36728 49292 36737
rect 52092 36771 52144 36780
rect 36728 36592 36780 36644
rect 42984 36660 43036 36712
rect 39488 36592 39540 36644
rect 38016 36524 38068 36576
rect 38384 36524 38436 36576
rect 39212 36524 39264 36576
rect 40592 36524 40644 36576
rect 42984 36524 43036 36576
rect 44180 36660 44232 36712
rect 46112 36660 46164 36712
rect 46848 36660 46900 36712
rect 49148 36703 49200 36712
rect 49148 36669 49157 36703
rect 49157 36669 49191 36703
rect 49191 36669 49200 36703
rect 49148 36660 49200 36669
rect 49700 36660 49752 36712
rect 48136 36635 48188 36644
rect 48136 36601 48145 36635
rect 48145 36601 48179 36635
rect 48179 36601 48188 36635
rect 48136 36592 48188 36601
rect 52092 36737 52101 36771
rect 52101 36737 52135 36771
rect 52135 36737 52144 36771
rect 52092 36728 52144 36737
rect 52276 36771 52328 36780
rect 52276 36737 52290 36771
rect 52290 36737 52324 36771
rect 52324 36737 52328 36771
rect 52276 36728 52328 36737
rect 53196 36771 53248 36780
rect 53196 36737 53205 36771
rect 53205 36737 53239 36771
rect 53239 36737 53248 36771
rect 53196 36728 53248 36737
rect 53472 36796 53524 36848
rect 53564 36771 53616 36780
rect 53564 36737 53573 36771
rect 53573 36737 53607 36771
rect 53607 36737 53616 36771
rect 53564 36728 53616 36737
rect 53656 36728 53708 36780
rect 54852 36703 54904 36712
rect 54852 36669 54861 36703
rect 54861 36669 54895 36703
rect 54895 36669 54904 36703
rect 54852 36660 54904 36669
rect 56232 36592 56284 36644
rect 43996 36524 44048 36576
rect 45100 36524 45152 36576
rect 46296 36524 46348 36576
rect 47400 36524 47452 36576
rect 47584 36524 47636 36576
rect 50068 36524 50120 36576
rect 50344 36567 50396 36576
rect 50344 36533 50353 36567
rect 50353 36533 50387 36567
rect 50387 36533 50396 36567
rect 50344 36524 50396 36533
rect 50712 36524 50764 36576
rect 52828 36524 52880 36576
rect 54208 36524 54260 36576
rect 54760 36524 54812 36576
rect 55128 36567 55180 36576
rect 55128 36533 55137 36567
rect 55137 36533 55171 36567
rect 55171 36533 55180 36567
rect 55128 36524 55180 36533
rect 56600 36524 56652 36576
rect 57980 36524 58032 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 29920 36320 29972 36372
rect 33140 36320 33192 36372
rect 34060 36320 34112 36372
rect 34244 36320 34296 36372
rect 36636 36320 36688 36372
rect 40224 36320 40276 36372
rect 41512 36320 41564 36372
rect 49240 36320 49292 36372
rect 29828 36295 29880 36304
rect 29828 36261 29837 36295
rect 29837 36261 29871 36295
rect 29871 36261 29880 36295
rect 29828 36252 29880 36261
rect 31484 36252 31536 36304
rect 33692 36252 33744 36304
rect 30380 36184 30432 36236
rect 30932 36227 30984 36236
rect 30932 36193 30941 36227
rect 30941 36193 30975 36227
rect 30975 36193 30984 36227
rect 30932 36184 30984 36193
rect 31392 36184 31444 36236
rect 28908 36159 28960 36168
rect 28908 36125 28917 36159
rect 28917 36125 28951 36159
rect 28951 36125 28960 36159
rect 28908 36116 28960 36125
rect 29276 36116 29328 36168
rect 30564 36159 30616 36168
rect 30564 36125 30573 36159
rect 30573 36125 30607 36159
rect 30607 36125 30616 36159
rect 30564 36116 30616 36125
rect 33048 36184 33100 36236
rect 33508 36159 33560 36168
rect 29184 36091 29236 36100
rect 29184 36057 29193 36091
rect 29193 36057 29227 36091
rect 29227 36057 29236 36091
rect 29184 36048 29236 36057
rect 29828 36048 29880 36100
rect 33508 36125 33517 36159
rect 33517 36125 33551 36159
rect 33551 36125 33560 36159
rect 33508 36116 33560 36125
rect 34060 36184 34112 36236
rect 33324 36048 33376 36100
rect 33784 36091 33836 36100
rect 33784 36057 33793 36091
rect 33793 36057 33827 36091
rect 33827 36057 33836 36091
rect 33784 36048 33836 36057
rect 28356 35980 28408 36032
rect 30656 35980 30708 36032
rect 32496 35980 32548 36032
rect 34888 36048 34940 36100
rect 35992 36116 36044 36168
rect 36728 36184 36780 36236
rect 37464 36184 37516 36236
rect 37188 36116 37240 36168
rect 37648 36159 37700 36168
rect 37648 36125 37657 36159
rect 37657 36125 37691 36159
rect 37691 36125 37700 36159
rect 37648 36116 37700 36125
rect 40592 36252 40644 36304
rect 42524 36252 42576 36304
rect 44916 36252 44968 36304
rect 46940 36252 46992 36304
rect 47952 36252 48004 36304
rect 39948 36184 40000 36236
rect 34060 35980 34112 36032
rect 34612 35980 34664 36032
rect 35900 35980 35952 36032
rect 36360 35980 36412 36032
rect 37556 36048 37608 36100
rect 38292 36116 38344 36168
rect 40132 36116 40184 36168
rect 41512 36184 41564 36236
rect 41788 36184 41840 36236
rect 42892 36227 42944 36236
rect 42892 36193 42901 36227
rect 42901 36193 42935 36227
rect 42935 36193 42944 36227
rect 42892 36184 42944 36193
rect 42984 36184 43036 36236
rect 45008 36184 45060 36236
rect 45744 36227 45796 36236
rect 45744 36193 45753 36227
rect 45753 36193 45787 36227
rect 45787 36193 45796 36227
rect 45744 36184 45796 36193
rect 41880 36159 41932 36168
rect 41880 36125 41889 36159
rect 41889 36125 41923 36159
rect 41923 36125 41932 36159
rect 41880 36116 41932 36125
rect 42340 36116 42392 36168
rect 38016 36091 38068 36100
rect 38016 36057 38025 36091
rect 38025 36057 38059 36091
rect 38059 36057 38068 36091
rect 38016 36048 38068 36057
rect 38384 35980 38436 36032
rect 42616 36116 42668 36168
rect 43168 36159 43220 36168
rect 43168 36125 43177 36159
rect 43177 36125 43211 36159
rect 43211 36125 43220 36159
rect 43168 36116 43220 36125
rect 38660 35980 38712 36032
rect 40132 35980 40184 36032
rect 40684 35980 40736 36032
rect 42708 35980 42760 36032
rect 44456 36159 44508 36168
rect 44456 36125 44465 36159
rect 44465 36125 44499 36159
rect 44499 36125 44508 36159
rect 44456 36116 44508 36125
rect 46480 36159 46532 36168
rect 46480 36125 46489 36159
rect 46489 36125 46523 36159
rect 46523 36125 46532 36159
rect 46480 36116 46532 36125
rect 44916 36048 44968 36100
rect 46848 36116 46900 36168
rect 47400 36159 47452 36168
rect 47400 36125 47409 36159
rect 47409 36125 47443 36159
rect 47443 36125 47452 36159
rect 47400 36116 47452 36125
rect 47584 36159 47636 36168
rect 47584 36125 47593 36159
rect 47593 36125 47627 36159
rect 47627 36125 47636 36159
rect 47584 36116 47636 36125
rect 48688 36184 48740 36236
rect 49700 36227 49752 36236
rect 49700 36193 49709 36227
rect 49709 36193 49743 36227
rect 49743 36193 49752 36227
rect 50712 36252 50764 36304
rect 49700 36184 49752 36193
rect 49056 36159 49108 36168
rect 49056 36125 49065 36159
rect 49065 36125 49099 36159
rect 49099 36125 49108 36159
rect 49056 36116 49108 36125
rect 50344 36159 50396 36168
rect 50344 36125 50353 36159
rect 50353 36125 50387 36159
rect 50387 36125 50396 36159
rect 50344 36116 50396 36125
rect 50988 36184 51040 36236
rect 52828 36227 52880 36236
rect 52828 36193 52837 36227
rect 52837 36193 52871 36227
rect 52871 36193 52880 36227
rect 52828 36184 52880 36193
rect 50620 36159 50672 36168
rect 50620 36125 50629 36159
rect 50629 36125 50663 36159
rect 50663 36125 50672 36159
rect 50620 36116 50672 36125
rect 50896 36116 50948 36168
rect 51264 36116 51316 36168
rect 52736 36159 52788 36168
rect 52736 36125 52745 36159
rect 52745 36125 52779 36159
rect 52779 36125 52788 36159
rect 52736 36116 52788 36125
rect 53288 36116 53340 36168
rect 53656 36116 53708 36168
rect 55128 36116 55180 36168
rect 56140 36159 56192 36168
rect 56140 36125 56149 36159
rect 56149 36125 56183 36159
rect 56183 36125 56192 36159
rect 56140 36116 56192 36125
rect 57428 36159 57480 36168
rect 57428 36125 57437 36159
rect 57437 36125 57471 36159
rect 57471 36125 57480 36159
rect 57428 36116 57480 36125
rect 57704 36159 57756 36168
rect 57704 36125 57713 36159
rect 57713 36125 57747 36159
rect 57747 36125 57756 36159
rect 57704 36116 57756 36125
rect 48412 36048 48464 36100
rect 50068 36048 50120 36100
rect 44272 35980 44324 36032
rect 45192 36023 45244 36032
rect 45192 35989 45201 36023
rect 45201 35989 45235 36023
rect 45235 35989 45244 36023
rect 45192 35980 45244 35989
rect 46572 36023 46624 36032
rect 46572 35989 46581 36023
rect 46581 35989 46615 36023
rect 46615 35989 46624 36023
rect 46572 35980 46624 35989
rect 47952 35980 48004 36032
rect 48136 36023 48188 36032
rect 48136 35989 48145 36023
rect 48145 35989 48179 36023
rect 48179 35989 48188 36023
rect 48136 35980 48188 35989
rect 48504 35980 48556 36032
rect 49332 35980 49384 36032
rect 50804 35980 50856 36032
rect 51632 36023 51684 36032
rect 51632 35989 51641 36023
rect 51641 35989 51675 36023
rect 51675 35989 51684 36023
rect 51632 35980 51684 35989
rect 52092 35980 52144 36032
rect 54300 35980 54352 36032
rect 54668 35980 54720 36032
rect 54852 36023 54904 36032
rect 54852 35989 54861 36023
rect 54861 35989 54895 36023
rect 54895 35989 54904 36023
rect 54852 35980 54904 35989
rect 55220 35980 55272 36032
rect 56876 35980 56928 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 29460 35776 29512 35828
rect 30288 35776 30340 35828
rect 31668 35776 31720 35828
rect 28908 35708 28960 35760
rect 29184 35640 29236 35692
rect 30104 35683 30156 35692
rect 30104 35649 30113 35683
rect 30113 35649 30147 35683
rect 30147 35649 30156 35683
rect 30104 35640 30156 35649
rect 30564 35708 30616 35760
rect 31300 35708 31352 35760
rect 31208 35683 31260 35692
rect 31208 35649 31217 35683
rect 31217 35649 31251 35683
rect 31251 35649 31260 35683
rect 31208 35640 31260 35649
rect 31392 35683 31444 35692
rect 31392 35649 31401 35683
rect 31401 35649 31435 35683
rect 31435 35649 31444 35683
rect 31392 35640 31444 35649
rect 33600 35751 33652 35760
rect 33600 35717 33609 35751
rect 33609 35717 33643 35751
rect 33643 35717 33652 35751
rect 33600 35708 33652 35717
rect 29276 35547 29328 35556
rect 29276 35513 29285 35547
rect 29285 35513 29319 35547
rect 29319 35513 29328 35547
rect 29276 35504 29328 35513
rect 33324 35640 33376 35692
rect 34060 35640 34112 35692
rect 34704 35776 34756 35828
rect 35716 35776 35768 35828
rect 34888 35708 34940 35760
rect 37464 35776 37516 35828
rect 38936 35776 38988 35828
rect 41420 35776 41472 35828
rect 42708 35819 42760 35828
rect 38844 35708 38896 35760
rect 42708 35785 42717 35819
rect 42717 35785 42751 35819
rect 42751 35785 42760 35819
rect 42708 35776 42760 35785
rect 43076 35819 43128 35828
rect 43076 35785 43085 35819
rect 43085 35785 43119 35819
rect 43119 35785 43128 35819
rect 43076 35776 43128 35785
rect 44456 35776 44508 35828
rect 32864 35615 32916 35624
rect 32864 35581 32873 35615
rect 32873 35581 32907 35615
rect 32907 35581 32916 35615
rect 32864 35572 32916 35581
rect 32772 35504 32824 35556
rect 32312 35479 32364 35488
rect 32312 35445 32321 35479
rect 32321 35445 32355 35479
rect 32355 35445 32364 35479
rect 32312 35436 32364 35445
rect 32404 35436 32456 35488
rect 32956 35504 33008 35556
rect 35348 35615 35400 35624
rect 35348 35581 35357 35615
rect 35357 35581 35391 35615
rect 35391 35581 35400 35615
rect 35348 35572 35400 35581
rect 35440 35504 35492 35556
rect 36544 35640 36596 35692
rect 37464 35683 37516 35692
rect 37464 35649 37473 35683
rect 37473 35649 37507 35683
rect 37507 35649 37516 35683
rect 37464 35640 37516 35649
rect 37556 35683 37608 35692
rect 37556 35649 37565 35683
rect 37565 35649 37599 35683
rect 37599 35649 37608 35683
rect 37556 35640 37608 35649
rect 37740 35683 37792 35692
rect 37740 35649 37749 35683
rect 37749 35649 37783 35683
rect 37783 35649 37792 35683
rect 38568 35683 38620 35692
rect 37740 35640 37792 35649
rect 38568 35649 38577 35683
rect 38577 35649 38611 35683
rect 38611 35649 38620 35683
rect 38568 35640 38620 35649
rect 39212 35683 39264 35692
rect 39212 35649 39221 35683
rect 39221 35649 39255 35683
rect 39255 35649 39264 35683
rect 39212 35640 39264 35649
rect 40868 35640 40920 35692
rect 41420 35683 41472 35692
rect 41420 35649 41429 35683
rect 41429 35649 41463 35683
rect 41463 35649 41472 35683
rect 41420 35640 41472 35649
rect 41880 35640 41932 35692
rect 42616 35683 42668 35692
rect 42616 35649 42625 35683
rect 42625 35649 42659 35683
rect 42659 35649 42668 35683
rect 42616 35640 42668 35649
rect 43168 35640 43220 35692
rect 44088 35683 44140 35692
rect 44088 35649 44097 35683
rect 44097 35649 44131 35683
rect 44131 35649 44140 35683
rect 44088 35640 44140 35649
rect 44180 35640 44232 35692
rect 45192 35683 45244 35692
rect 45192 35649 45201 35683
rect 45201 35649 45235 35683
rect 45235 35649 45244 35683
rect 45192 35640 45244 35649
rect 45744 35776 45796 35828
rect 46112 35708 46164 35760
rect 45928 35640 45980 35692
rect 46204 35683 46256 35692
rect 46204 35649 46213 35683
rect 46213 35649 46247 35683
rect 46247 35649 46256 35683
rect 46204 35640 46256 35649
rect 47952 35683 48004 35692
rect 37188 35504 37240 35556
rect 37648 35504 37700 35556
rect 47952 35649 47961 35683
rect 47961 35649 47995 35683
rect 47995 35649 48004 35683
rect 47952 35640 48004 35649
rect 40960 35504 41012 35556
rect 36176 35436 36228 35488
rect 47124 35572 47176 35624
rect 47308 35572 47360 35624
rect 50620 35751 50672 35760
rect 48780 35683 48832 35692
rect 48780 35649 48789 35683
rect 48789 35649 48823 35683
rect 48823 35649 48832 35683
rect 48780 35640 48832 35649
rect 48872 35572 48924 35624
rect 44088 35504 44140 35556
rect 46204 35504 46256 35556
rect 48320 35547 48372 35556
rect 48320 35513 48329 35547
rect 48329 35513 48363 35547
rect 48363 35513 48372 35547
rect 48320 35504 48372 35513
rect 48688 35504 48740 35556
rect 50252 35640 50304 35692
rect 50620 35717 50629 35751
rect 50629 35717 50663 35751
rect 50663 35717 50672 35751
rect 50620 35708 50672 35717
rect 50988 35776 51040 35828
rect 52276 35776 52328 35828
rect 50712 35683 50764 35692
rect 49976 35504 50028 35556
rect 45468 35436 45520 35488
rect 46664 35479 46716 35488
rect 46664 35445 46673 35479
rect 46673 35445 46707 35479
rect 46707 35445 46716 35479
rect 46664 35436 46716 35445
rect 50712 35649 50721 35683
rect 50721 35649 50755 35683
rect 50755 35649 50764 35683
rect 50712 35640 50764 35649
rect 54668 35708 54720 35760
rect 50620 35572 50672 35624
rect 52736 35640 52788 35692
rect 53656 35640 53708 35692
rect 54576 35683 54628 35692
rect 54576 35649 54586 35683
rect 54586 35649 54620 35683
rect 54620 35649 54628 35683
rect 57428 35776 57480 35828
rect 56692 35708 56744 35760
rect 57336 35751 57388 35760
rect 57336 35717 57345 35751
rect 57345 35717 57379 35751
rect 57379 35717 57388 35751
rect 57336 35708 57388 35717
rect 54576 35640 54628 35649
rect 50896 35504 50948 35556
rect 53472 35572 53524 35624
rect 51908 35436 51960 35488
rect 56140 35640 56192 35692
rect 54760 35572 54812 35624
rect 55404 35436 55456 35488
rect 57704 35436 57756 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 30104 35232 30156 35284
rect 31208 35232 31260 35284
rect 32036 35232 32088 35284
rect 32772 35207 32824 35216
rect 32772 35173 32781 35207
rect 32781 35173 32815 35207
rect 32815 35173 32824 35207
rect 32772 35164 32824 35173
rect 33508 35232 33560 35284
rect 33876 35232 33928 35284
rect 35440 35275 35492 35284
rect 35440 35241 35449 35275
rect 35449 35241 35483 35275
rect 35483 35241 35492 35275
rect 35440 35232 35492 35241
rect 33968 35164 34020 35216
rect 37740 35232 37792 35284
rect 37832 35232 37884 35284
rect 41972 35232 42024 35284
rect 47308 35275 47360 35284
rect 28908 35096 28960 35148
rect 29000 35071 29052 35080
rect 29000 35037 29009 35071
rect 29009 35037 29043 35071
rect 29043 35037 29052 35071
rect 29000 35028 29052 35037
rect 30656 35071 30708 35080
rect 27344 34960 27396 35012
rect 30656 35037 30665 35071
rect 30665 35037 30699 35071
rect 30699 35037 30708 35071
rect 30656 35028 30708 35037
rect 31300 35071 31352 35080
rect 31300 35037 31309 35071
rect 31309 35037 31343 35071
rect 31343 35037 31352 35071
rect 31300 35028 31352 35037
rect 31760 35028 31812 35080
rect 32404 35071 32456 35080
rect 32404 35037 32413 35071
rect 32413 35037 32447 35071
rect 32447 35037 32456 35071
rect 32404 35028 32456 35037
rect 31208 34960 31260 35012
rect 32036 34960 32088 35012
rect 32772 35071 32824 35080
rect 32772 35037 32781 35071
rect 32781 35037 32815 35071
rect 32815 35037 32824 35071
rect 32772 35028 32824 35037
rect 33324 35028 33376 35080
rect 33692 35071 33744 35080
rect 33692 35037 33701 35071
rect 33701 35037 33735 35071
rect 33735 35037 33744 35071
rect 33692 35028 33744 35037
rect 33784 34960 33836 35012
rect 35716 35028 35768 35080
rect 36176 35096 36228 35148
rect 38200 35164 38252 35216
rect 38660 35164 38712 35216
rect 47308 35241 47317 35275
rect 47317 35241 47351 35275
rect 47351 35241 47360 35275
rect 47308 35232 47360 35241
rect 49700 35275 49752 35284
rect 49700 35241 49709 35275
rect 49709 35241 49743 35275
rect 49743 35241 49752 35275
rect 49700 35232 49752 35241
rect 52552 35232 52604 35284
rect 53656 35275 53708 35284
rect 53656 35241 53665 35275
rect 53665 35241 53699 35275
rect 53699 35241 53708 35275
rect 53656 35232 53708 35241
rect 37188 35139 37240 35148
rect 37188 35105 37197 35139
rect 37197 35105 37231 35139
rect 37231 35105 37240 35139
rect 37188 35096 37240 35105
rect 36176 34960 36228 35012
rect 37004 35071 37056 35080
rect 37004 35037 37013 35071
rect 37013 35037 37047 35071
rect 37047 35037 37056 35071
rect 37464 35096 37516 35148
rect 43260 35096 43312 35148
rect 43536 35164 43588 35216
rect 49056 35164 49108 35216
rect 37004 35028 37056 35037
rect 37740 35028 37792 35080
rect 38200 35071 38252 35080
rect 38200 35037 38209 35071
rect 38209 35037 38243 35071
rect 38243 35037 38252 35071
rect 38200 35028 38252 35037
rect 37648 34960 37700 35012
rect 38936 35028 38988 35080
rect 41144 35028 41196 35080
rect 41420 35028 41472 35080
rect 41880 35071 41932 35080
rect 40132 35003 40184 35012
rect 40132 34969 40141 35003
rect 40141 34969 40175 35003
rect 40175 34969 40184 35003
rect 40132 34960 40184 34969
rect 41512 34960 41564 35012
rect 41880 35037 41889 35071
rect 41889 35037 41923 35071
rect 41923 35037 41932 35071
rect 41880 35028 41932 35037
rect 43168 35028 43220 35080
rect 43996 35071 44048 35080
rect 43996 35037 44005 35071
rect 44005 35037 44039 35071
rect 44039 35037 44048 35071
rect 43996 35028 44048 35037
rect 42340 34960 42392 35012
rect 42984 34960 43036 35012
rect 30472 34892 30524 34944
rect 32680 34892 32732 34944
rect 34520 34892 34572 34944
rect 35440 34892 35492 34944
rect 35808 34935 35860 34944
rect 35808 34901 35817 34935
rect 35817 34901 35851 34935
rect 35851 34901 35860 34935
rect 35808 34892 35860 34901
rect 37556 34892 37608 34944
rect 38844 34892 38896 34944
rect 41696 34892 41748 34944
rect 42524 34892 42576 34944
rect 45928 35096 45980 35148
rect 46664 35071 46716 35080
rect 46664 35037 46673 35071
rect 46673 35037 46707 35071
rect 46707 35037 46716 35071
rect 46664 35028 46716 35037
rect 47860 35096 47912 35148
rect 46940 35071 46992 35080
rect 46940 35037 46949 35071
rect 46949 35037 46983 35071
rect 46983 35037 46992 35071
rect 46940 35028 46992 35037
rect 48136 35028 48188 35080
rect 48320 35096 48372 35148
rect 53748 35164 53800 35216
rect 55772 35164 55824 35216
rect 56600 35164 56652 35216
rect 58072 35164 58124 35216
rect 48688 35028 48740 35080
rect 48872 35071 48924 35080
rect 48872 35037 48881 35071
rect 48881 35037 48915 35071
rect 48915 35037 48924 35071
rect 48872 35028 48924 35037
rect 50804 35071 50856 35080
rect 47584 34960 47636 35012
rect 48320 34960 48372 35012
rect 48780 34960 48832 35012
rect 50804 35037 50813 35071
rect 50813 35037 50847 35071
rect 50847 35037 50856 35071
rect 50804 35028 50856 35037
rect 53196 35028 53248 35080
rect 49976 34960 50028 35012
rect 53380 34960 53432 35012
rect 54760 35028 54812 35080
rect 55496 35096 55548 35148
rect 57980 35096 58032 35148
rect 55772 35028 55824 35080
rect 56140 35071 56192 35080
rect 56140 35037 56149 35071
rect 56149 35037 56183 35071
rect 56183 35037 56192 35071
rect 56140 35028 56192 35037
rect 56324 35028 56376 35080
rect 57152 35071 57204 35080
rect 57152 35037 57161 35071
rect 57161 35037 57195 35071
rect 57195 35037 57204 35071
rect 57152 35028 57204 35037
rect 57336 35071 57388 35080
rect 57336 35037 57345 35071
rect 57345 35037 57379 35071
rect 57379 35037 57388 35071
rect 57336 35028 57388 35037
rect 57704 34960 57756 35012
rect 43904 34935 43956 34944
rect 43904 34901 43913 34935
rect 43913 34901 43947 34935
rect 43947 34901 43956 34935
rect 43904 34892 43956 34901
rect 44456 34935 44508 34944
rect 44456 34901 44465 34935
rect 44465 34901 44499 34935
rect 44499 34901 44508 34935
rect 44456 34892 44508 34901
rect 45192 34892 45244 34944
rect 46940 34892 46992 34944
rect 47952 34892 48004 34944
rect 51356 34892 51408 34944
rect 52644 34892 52696 34944
rect 54116 34892 54168 34944
rect 55956 34892 56008 34944
rect 56968 34935 57020 34944
rect 56968 34901 56977 34935
rect 56977 34901 57011 34935
rect 57011 34901 57020 34935
rect 56968 34892 57020 34901
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 27620 34688 27672 34740
rect 29000 34688 29052 34740
rect 32496 34731 32548 34740
rect 29092 34620 29144 34672
rect 30196 34620 30248 34672
rect 30656 34620 30708 34672
rect 27344 34595 27396 34604
rect 27344 34561 27353 34595
rect 27353 34561 27387 34595
rect 27387 34561 27396 34595
rect 27344 34552 27396 34561
rect 31208 34552 31260 34604
rect 31760 34620 31812 34672
rect 28080 34527 28132 34536
rect 28080 34493 28089 34527
rect 28089 34493 28123 34527
rect 28123 34493 28132 34527
rect 28080 34484 28132 34493
rect 31668 34484 31720 34536
rect 32496 34697 32505 34731
rect 32505 34697 32539 34731
rect 32539 34697 32548 34731
rect 32496 34688 32548 34697
rect 32680 34688 32732 34740
rect 31944 34620 31996 34672
rect 33232 34620 33284 34672
rect 35348 34620 35400 34672
rect 37004 34620 37056 34672
rect 33140 34595 33192 34604
rect 33140 34561 33149 34595
rect 33149 34561 33183 34595
rect 33183 34561 33192 34595
rect 33140 34552 33192 34561
rect 33784 34595 33836 34604
rect 33784 34561 33793 34595
rect 33793 34561 33827 34595
rect 33827 34561 33836 34595
rect 33784 34552 33836 34561
rect 34336 34484 34388 34536
rect 35348 34484 35400 34536
rect 35532 34595 35584 34604
rect 35532 34561 35541 34595
rect 35541 34561 35575 34595
rect 35575 34561 35584 34595
rect 35532 34552 35584 34561
rect 38660 34620 38712 34672
rect 39304 34620 39356 34672
rect 40316 34663 40368 34672
rect 40316 34629 40325 34663
rect 40325 34629 40359 34663
rect 40359 34629 40368 34663
rect 40316 34620 40368 34629
rect 41052 34688 41104 34740
rect 42340 34688 42392 34740
rect 43720 34688 43772 34740
rect 44456 34688 44508 34740
rect 48964 34688 49016 34740
rect 50988 34688 51040 34740
rect 33416 34416 33468 34468
rect 28540 34348 28592 34400
rect 32312 34348 32364 34400
rect 32772 34348 32824 34400
rect 33048 34348 33100 34400
rect 37188 34484 37240 34536
rect 37648 34552 37700 34604
rect 38292 34595 38344 34604
rect 38292 34561 38301 34595
rect 38301 34561 38335 34595
rect 38335 34561 38344 34595
rect 38292 34552 38344 34561
rect 41972 34552 42024 34604
rect 43168 34552 43220 34604
rect 44088 34552 44140 34604
rect 45928 34620 45980 34672
rect 45836 34552 45888 34604
rect 46112 34552 46164 34604
rect 46572 34552 46624 34604
rect 37832 34484 37884 34536
rect 41052 34527 41104 34536
rect 41052 34493 41061 34527
rect 41061 34493 41095 34527
rect 41095 34493 41104 34527
rect 41052 34484 41104 34493
rect 41144 34484 41196 34536
rect 43536 34527 43588 34536
rect 43536 34493 43545 34527
rect 43545 34493 43579 34527
rect 43579 34493 43588 34527
rect 43536 34484 43588 34493
rect 45100 34527 45152 34536
rect 45100 34493 45109 34527
rect 45109 34493 45143 34527
rect 45143 34493 45152 34527
rect 45100 34484 45152 34493
rect 36176 34391 36228 34400
rect 36176 34357 36185 34391
rect 36185 34357 36219 34391
rect 36219 34357 36228 34391
rect 36176 34348 36228 34357
rect 37648 34391 37700 34400
rect 37648 34357 37657 34391
rect 37657 34357 37691 34391
rect 37691 34357 37700 34391
rect 37648 34348 37700 34357
rect 39120 34348 39172 34400
rect 44180 34348 44232 34400
rect 44548 34348 44600 34400
rect 48872 34620 48924 34672
rect 49608 34620 49660 34672
rect 52368 34620 52420 34672
rect 47860 34552 47912 34604
rect 48320 34552 48372 34604
rect 48688 34552 48740 34604
rect 49332 34595 49384 34604
rect 49332 34561 49341 34595
rect 49341 34561 49375 34595
rect 49375 34561 49384 34595
rect 49332 34552 49384 34561
rect 50804 34552 50856 34604
rect 51448 34552 51500 34604
rect 51724 34595 51776 34604
rect 51724 34561 51733 34595
rect 51733 34561 51767 34595
rect 51767 34561 51776 34595
rect 51724 34552 51776 34561
rect 52920 34595 52972 34604
rect 52920 34561 52929 34595
rect 52929 34561 52963 34595
rect 52963 34561 52972 34595
rect 52920 34552 52972 34561
rect 56324 34688 56376 34740
rect 57152 34688 57204 34740
rect 54576 34620 54628 34672
rect 55496 34595 55548 34604
rect 55496 34561 55505 34595
rect 55505 34561 55539 34595
rect 55539 34561 55548 34595
rect 55496 34552 55548 34561
rect 56324 34595 56376 34604
rect 56324 34561 56333 34595
rect 56333 34561 56367 34595
rect 56367 34561 56376 34595
rect 56324 34552 56376 34561
rect 57980 34620 58032 34672
rect 58072 34595 58124 34604
rect 51540 34484 51592 34536
rect 55588 34527 55640 34536
rect 55588 34493 55597 34527
rect 55597 34493 55631 34527
rect 55631 34493 55640 34527
rect 55588 34484 55640 34493
rect 56140 34484 56192 34536
rect 58072 34561 58081 34595
rect 58081 34561 58115 34595
rect 58115 34561 58124 34595
rect 58072 34552 58124 34561
rect 57060 34527 57112 34536
rect 57060 34493 57069 34527
rect 57069 34493 57103 34527
rect 57103 34493 57112 34527
rect 57060 34484 57112 34493
rect 52460 34416 52512 34468
rect 52920 34416 52972 34468
rect 46296 34391 46348 34400
rect 46296 34357 46305 34391
rect 46305 34357 46339 34391
rect 46339 34357 46348 34391
rect 46296 34348 46348 34357
rect 47860 34391 47912 34400
rect 47860 34357 47869 34391
rect 47869 34357 47903 34391
rect 47903 34357 47912 34391
rect 47860 34348 47912 34357
rect 49976 34348 50028 34400
rect 53380 34348 53432 34400
rect 54484 34348 54536 34400
rect 56048 34348 56100 34400
rect 57336 34348 57388 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 28080 34144 28132 34196
rect 29092 34187 29144 34196
rect 29092 34153 29101 34187
rect 29101 34153 29135 34187
rect 29135 34153 29144 34187
rect 29092 34144 29144 34153
rect 30656 34144 30708 34196
rect 33140 34144 33192 34196
rect 36360 34144 36412 34196
rect 37372 34144 37424 34196
rect 39304 34144 39356 34196
rect 43260 34187 43312 34196
rect 43260 34153 43269 34187
rect 43269 34153 43303 34187
rect 43303 34153 43312 34187
rect 43260 34144 43312 34153
rect 43904 34144 43956 34196
rect 45836 34144 45888 34196
rect 48596 34144 48648 34196
rect 52092 34144 52144 34196
rect 57704 34187 57756 34196
rect 57704 34153 57713 34187
rect 57713 34153 57747 34187
rect 57747 34153 57756 34187
rect 57704 34144 57756 34153
rect 45560 34076 45612 34128
rect 29736 34008 29788 34060
rect 29184 33940 29236 33992
rect 31668 33940 31720 33992
rect 27620 33915 27672 33924
rect 27620 33881 27629 33915
rect 27629 33881 27663 33915
rect 27663 33881 27672 33915
rect 27620 33872 27672 33881
rect 28908 33872 28960 33924
rect 30564 33872 30616 33924
rect 34336 34008 34388 34060
rect 33048 33940 33100 33992
rect 33324 33872 33376 33924
rect 33600 33983 33652 33992
rect 33600 33949 33609 33983
rect 33609 33949 33643 33983
rect 33643 33949 33652 33983
rect 33600 33940 33652 33949
rect 33784 33983 33836 33992
rect 33784 33949 33793 33983
rect 33793 33949 33827 33983
rect 33827 33949 33836 33983
rect 33784 33940 33836 33949
rect 36544 34008 36596 34060
rect 37556 34008 37608 34060
rect 38660 34008 38712 34060
rect 40224 34008 40276 34060
rect 41696 34008 41748 34060
rect 42340 34051 42392 34060
rect 42340 34017 42349 34051
rect 42349 34017 42383 34051
rect 42383 34017 42392 34051
rect 42340 34008 42392 34017
rect 42984 34008 43036 34060
rect 43628 34008 43680 34060
rect 44180 34051 44232 34060
rect 44180 34017 44189 34051
rect 44189 34017 44223 34051
rect 44223 34017 44232 34051
rect 44180 34008 44232 34017
rect 36176 33872 36228 33924
rect 37648 33872 37700 33924
rect 37832 33872 37884 33924
rect 38016 33872 38068 33924
rect 38844 33872 38896 33924
rect 37096 33847 37148 33856
rect 37096 33813 37105 33847
rect 37105 33813 37139 33847
rect 37139 33813 37148 33847
rect 37096 33804 37148 33813
rect 43168 33940 43220 33992
rect 43352 33940 43404 33992
rect 50620 34076 50672 34128
rect 51632 34076 51684 34128
rect 54208 34119 54260 34128
rect 46388 34008 46440 34060
rect 49976 34008 50028 34060
rect 45836 33983 45888 33992
rect 45836 33949 45845 33983
rect 45845 33949 45879 33983
rect 45879 33949 45888 33983
rect 45836 33940 45888 33949
rect 41972 33872 42024 33924
rect 42064 33872 42116 33924
rect 42616 33872 42668 33924
rect 42800 33804 42852 33856
rect 43260 33804 43312 33856
rect 46204 33847 46256 33856
rect 46204 33813 46213 33847
rect 46213 33813 46247 33847
rect 46247 33813 46256 33847
rect 46204 33804 46256 33813
rect 48688 33983 48740 33992
rect 48688 33949 48697 33983
rect 48697 33949 48731 33983
rect 48731 33949 48740 33983
rect 48688 33940 48740 33949
rect 48780 33940 48832 33992
rect 49608 33983 49660 33992
rect 49608 33949 49617 33983
rect 49617 33949 49651 33983
rect 49651 33949 49660 33983
rect 49608 33940 49660 33949
rect 50988 33983 51040 33992
rect 50988 33949 50997 33983
rect 50997 33949 51031 33983
rect 51031 33949 51040 33983
rect 50988 33940 51040 33949
rect 52092 33983 52144 33992
rect 47768 33872 47820 33924
rect 48596 33872 48648 33924
rect 49332 33872 49384 33924
rect 49700 33872 49752 33924
rect 52092 33949 52101 33983
rect 52101 33949 52135 33983
rect 52135 33949 52144 33983
rect 52092 33940 52144 33949
rect 48320 33804 48372 33856
rect 50252 33804 50304 33856
rect 51356 33872 51408 33924
rect 51632 33804 51684 33856
rect 52000 33847 52052 33856
rect 52000 33813 52009 33847
rect 52009 33813 52043 33847
rect 52043 33813 52052 33847
rect 52000 33804 52052 33813
rect 53012 33847 53064 33856
rect 53012 33813 53021 33847
rect 53021 33813 53055 33847
rect 53055 33813 53064 33847
rect 53012 33804 53064 33813
rect 54208 34085 54217 34119
rect 54217 34085 54251 34119
rect 54251 34085 54260 34119
rect 54208 34076 54260 34085
rect 54024 33940 54076 33992
rect 54484 33983 54536 33992
rect 54484 33949 54493 33983
rect 54493 33949 54527 33983
rect 54527 33949 54536 33983
rect 54484 33940 54536 33949
rect 55956 33983 56008 33992
rect 55956 33949 55965 33983
rect 55965 33949 55999 33983
rect 55999 33949 56008 33983
rect 55956 33940 56008 33949
rect 56048 33983 56100 33992
rect 56048 33949 56057 33983
rect 56057 33949 56091 33983
rect 56091 33949 56100 33983
rect 56232 33983 56284 33992
rect 56048 33940 56100 33949
rect 56232 33949 56241 33983
rect 56241 33949 56275 33983
rect 56275 33949 56284 33983
rect 56232 33940 56284 33949
rect 56968 33940 57020 33992
rect 53564 33872 53616 33924
rect 55772 33872 55824 33924
rect 55864 33872 55916 33924
rect 56600 33872 56652 33924
rect 54392 33847 54444 33856
rect 54392 33813 54401 33847
rect 54401 33813 54435 33847
rect 54435 33813 54444 33847
rect 54392 33804 54444 33813
rect 56784 33847 56836 33856
rect 56784 33813 56793 33847
rect 56793 33813 56827 33847
rect 56827 33813 56836 33847
rect 56784 33804 56836 33813
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 31024 33532 31076 33584
rect 33600 33600 33652 33652
rect 34704 33600 34756 33652
rect 38844 33600 38896 33652
rect 41972 33643 42024 33652
rect 31760 33532 31812 33584
rect 33784 33532 33836 33584
rect 28080 33464 28132 33516
rect 29736 33507 29788 33516
rect 29736 33473 29745 33507
rect 29745 33473 29779 33507
rect 29779 33473 29788 33507
rect 29736 33464 29788 33473
rect 33232 33507 33284 33516
rect 33232 33473 33241 33507
rect 33241 33473 33275 33507
rect 33275 33473 33284 33507
rect 33232 33464 33284 33473
rect 34704 33507 34756 33516
rect 29184 33303 29236 33312
rect 29184 33269 29193 33303
rect 29193 33269 29227 33303
rect 29227 33269 29236 33303
rect 29184 33260 29236 33269
rect 33048 33396 33100 33448
rect 34704 33473 34713 33507
rect 34713 33473 34747 33507
rect 34747 33473 34756 33507
rect 38936 33532 38988 33584
rect 41972 33609 41981 33643
rect 41981 33609 42015 33643
rect 42015 33609 42024 33643
rect 41972 33600 42024 33609
rect 47216 33600 47268 33652
rect 49700 33600 49752 33652
rect 53564 33643 53616 33652
rect 34704 33464 34756 33473
rect 37280 33464 37332 33516
rect 37740 33464 37792 33516
rect 39488 33464 39540 33516
rect 42064 33507 42116 33516
rect 42064 33473 42073 33507
rect 42073 33473 42107 33507
rect 42107 33473 42116 33507
rect 42064 33464 42116 33473
rect 43352 33464 43404 33516
rect 45468 33532 45520 33584
rect 43904 33464 43956 33516
rect 44548 33507 44600 33516
rect 44548 33473 44557 33507
rect 44557 33473 44591 33507
rect 44591 33473 44600 33507
rect 44548 33464 44600 33473
rect 44640 33507 44692 33516
rect 44640 33473 44649 33507
rect 44649 33473 44683 33507
rect 44683 33473 44692 33507
rect 44640 33464 44692 33473
rect 46020 33507 46072 33516
rect 37096 33396 37148 33448
rect 38200 33439 38252 33448
rect 34612 33260 34664 33312
rect 35440 33328 35492 33380
rect 38200 33405 38209 33439
rect 38209 33405 38243 33439
rect 38243 33405 38252 33439
rect 38200 33396 38252 33405
rect 42708 33439 42760 33448
rect 42708 33405 42717 33439
rect 42717 33405 42751 33439
rect 42751 33405 42760 33439
rect 42708 33396 42760 33405
rect 43168 33396 43220 33448
rect 46020 33473 46029 33507
rect 46029 33473 46063 33507
rect 46063 33473 46072 33507
rect 46020 33464 46072 33473
rect 48228 33507 48280 33516
rect 48228 33473 48237 33507
rect 48237 33473 48271 33507
rect 48271 33473 48280 33507
rect 48228 33464 48280 33473
rect 48504 33507 48556 33516
rect 48504 33473 48513 33507
rect 48513 33473 48547 33507
rect 48547 33473 48556 33507
rect 48504 33464 48556 33473
rect 48688 33507 48740 33516
rect 48688 33473 48697 33507
rect 48697 33473 48731 33507
rect 48731 33473 48740 33507
rect 48688 33464 48740 33473
rect 49976 33507 50028 33516
rect 49976 33473 49985 33507
rect 49985 33473 50019 33507
rect 50019 33473 50028 33507
rect 49976 33464 50028 33473
rect 50252 33507 50304 33516
rect 50252 33473 50261 33507
rect 50261 33473 50295 33507
rect 50295 33473 50304 33507
rect 50252 33464 50304 33473
rect 52000 33532 52052 33584
rect 51356 33507 51408 33516
rect 51356 33473 51365 33507
rect 51365 33473 51399 33507
rect 51399 33473 51408 33507
rect 51356 33464 51408 33473
rect 52460 33532 52512 33584
rect 53564 33609 53573 33643
rect 53573 33609 53607 33643
rect 53607 33609 53616 33643
rect 53564 33600 53616 33609
rect 54024 33643 54076 33652
rect 54024 33609 54033 33643
rect 54033 33609 54067 33643
rect 54067 33609 54076 33643
rect 54024 33600 54076 33609
rect 57060 33600 57112 33652
rect 57428 33643 57480 33652
rect 57428 33609 57437 33643
rect 57437 33609 57471 33643
rect 57471 33609 57480 33643
rect 57428 33600 57480 33609
rect 53656 33532 53708 33584
rect 52368 33507 52420 33516
rect 52368 33473 52377 33507
rect 52377 33473 52411 33507
rect 52411 33473 52420 33507
rect 52368 33464 52420 33473
rect 53196 33507 53248 33516
rect 48412 33439 48464 33448
rect 48412 33405 48421 33439
rect 48421 33405 48455 33439
rect 48455 33405 48464 33439
rect 48412 33396 48464 33405
rect 49792 33396 49844 33448
rect 50988 33439 51040 33448
rect 50988 33405 50997 33439
rect 50997 33405 51031 33439
rect 51031 33405 51040 33439
rect 50988 33396 51040 33405
rect 51080 33396 51132 33448
rect 53196 33473 53205 33507
rect 53205 33473 53239 33507
rect 53239 33473 53248 33507
rect 53196 33464 53248 33473
rect 53380 33507 53432 33516
rect 53380 33473 53389 33507
rect 53389 33473 53423 33507
rect 53423 33473 53432 33507
rect 53380 33464 53432 33473
rect 54208 33507 54260 33516
rect 54208 33473 54217 33507
rect 54217 33473 54251 33507
rect 54251 33473 54260 33507
rect 54208 33464 54260 33473
rect 54484 33532 54536 33584
rect 56600 33464 56652 33516
rect 57520 33507 57572 33516
rect 57520 33473 57529 33507
rect 57529 33473 57563 33507
rect 57563 33473 57572 33507
rect 57520 33464 57572 33473
rect 53104 33439 53156 33448
rect 36728 33260 36780 33312
rect 37096 33260 37148 33312
rect 42984 33328 43036 33380
rect 46388 33328 46440 33380
rect 47860 33328 47912 33380
rect 50068 33371 50120 33380
rect 50068 33337 50077 33371
rect 50077 33337 50111 33371
rect 50111 33337 50120 33371
rect 50068 33328 50120 33337
rect 53104 33405 53113 33439
rect 53113 33405 53147 33439
rect 53147 33405 53156 33439
rect 53104 33396 53156 33405
rect 54484 33439 54536 33448
rect 38292 33260 38344 33312
rect 41420 33260 41472 33312
rect 41512 33260 41564 33312
rect 45192 33260 45244 33312
rect 45928 33260 45980 33312
rect 47032 33260 47084 33312
rect 49608 33260 49660 33312
rect 49700 33260 49752 33312
rect 49976 33260 50028 33312
rect 54484 33405 54493 33439
rect 54493 33405 54527 33439
rect 54527 33405 54536 33439
rect 54484 33396 54536 33405
rect 54944 33396 54996 33448
rect 56784 33396 56836 33448
rect 57888 33396 57940 33448
rect 57980 33396 58032 33448
rect 54116 33328 54168 33380
rect 55404 33328 55456 33380
rect 56692 33328 56744 33380
rect 53656 33260 53708 33312
rect 57980 33260 58032 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 29184 33099 29236 33108
rect 29184 33065 29193 33099
rect 29193 33065 29227 33099
rect 29227 33065 29236 33099
rect 29184 33056 29236 33065
rect 30564 33099 30616 33108
rect 30564 33065 30573 33099
rect 30573 33065 30607 33099
rect 30607 33065 30616 33099
rect 30564 33056 30616 33065
rect 34152 33056 34204 33108
rect 34612 33056 34664 33108
rect 35348 33056 35400 33108
rect 36544 33099 36596 33108
rect 29736 32920 29788 32972
rect 29184 32852 29236 32904
rect 30288 32852 30340 32904
rect 32864 32852 32916 32904
rect 34796 32852 34848 32904
rect 36544 33065 36553 33099
rect 36553 33065 36587 33099
rect 36587 33065 36596 33099
rect 36544 33056 36596 33065
rect 38936 33056 38988 33108
rect 41880 33099 41932 33108
rect 36728 32988 36780 33040
rect 36912 32920 36964 32972
rect 31576 32827 31628 32836
rect 31576 32793 31585 32827
rect 31585 32793 31619 32827
rect 31619 32793 31628 32827
rect 31576 32784 31628 32793
rect 37188 32852 37240 32904
rect 37372 32895 37424 32904
rect 37372 32861 37381 32895
rect 37381 32861 37415 32895
rect 37415 32861 37424 32895
rect 37372 32852 37424 32861
rect 39856 32920 39908 32972
rect 41052 32920 41104 32972
rect 41880 33065 41889 33099
rect 41889 33065 41923 33099
rect 41923 33065 41932 33099
rect 41880 33056 41932 33065
rect 48412 33056 48464 33108
rect 49792 33099 49844 33108
rect 49792 33065 49801 33099
rect 49801 33065 49835 33099
rect 49835 33065 49844 33099
rect 49792 33056 49844 33065
rect 50068 33056 50120 33108
rect 50804 33056 50856 33108
rect 37740 32895 37792 32904
rect 37740 32861 37749 32895
rect 37749 32861 37783 32895
rect 37783 32861 37792 32895
rect 37740 32852 37792 32861
rect 37924 32852 37976 32904
rect 38568 32852 38620 32904
rect 38660 32852 38712 32904
rect 39488 32852 39540 32904
rect 42340 32852 42392 32904
rect 42708 32852 42760 32904
rect 44640 32920 44692 32972
rect 46204 32963 46256 32972
rect 29644 32716 29696 32768
rect 37280 32784 37332 32836
rect 37648 32784 37700 32836
rect 40408 32827 40460 32836
rect 35992 32716 36044 32768
rect 38660 32716 38712 32768
rect 40408 32793 40417 32827
rect 40417 32793 40451 32827
rect 40451 32793 40460 32827
rect 40408 32784 40460 32793
rect 41420 32784 41472 32836
rect 40592 32716 40644 32768
rect 42800 32716 42852 32768
rect 43352 32852 43404 32904
rect 44088 32852 44140 32904
rect 46204 32929 46213 32963
rect 46213 32929 46247 32963
rect 46247 32929 46256 32963
rect 46204 32920 46256 32929
rect 48780 32988 48832 33040
rect 47584 32920 47636 32972
rect 43076 32784 43128 32836
rect 43536 32784 43588 32836
rect 46848 32852 46900 32904
rect 47400 32895 47452 32904
rect 47400 32861 47409 32895
rect 47409 32861 47443 32895
rect 47443 32861 47452 32895
rect 47400 32852 47452 32861
rect 48596 32852 48648 32904
rect 48412 32784 48464 32836
rect 51080 32920 51132 32972
rect 49608 32895 49660 32904
rect 49608 32861 49617 32895
rect 49617 32861 49651 32895
rect 49651 32861 49660 32895
rect 49608 32852 49660 32861
rect 49792 32895 49844 32904
rect 49792 32861 49801 32895
rect 49801 32861 49835 32895
rect 49835 32861 49844 32895
rect 52368 33056 52420 33108
rect 54576 33056 54628 33108
rect 55588 33056 55640 33108
rect 55772 32988 55824 33040
rect 56692 33056 56744 33108
rect 57520 33099 57572 33108
rect 57520 33065 57529 33099
rect 57529 33065 57563 33099
rect 57563 33065 57572 33099
rect 57520 33056 57572 33065
rect 52276 32920 52328 32972
rect 49792 32852 49844 32861
rect 50712 32784 50764 32836
rect 51632 32784 51684 32836
rect 52552 32895 52604 32904
rect 52552 32861 52561 32895
rect 52561 32861 52595 32895
rect 52595 32861 52604 32895
rect 52552 32852 52604 32861
rect 52920 32852 52972 32904
rect 53932 32895 53984 32904
rect 53932 32861 53941 32895
rect 53941 32861 53975 32895
rect 53975 32861 53984 32895
rect 53932 32852 53984 32861
rect 54116 32852 54168 32904
rect 54300 32895 54352 32904
rect 54300 32861 54309 32895
rect 54309 32861 54343 32895
rect 54343 32861 54352 32895
rect 54300 32852 54352 32861
rect 53564 32784 53616 32836
rect 55772 32895 55824 32904
rect 55772 32861 55781 32895
rect 55781 32861 55815 32895
rect 55815 32861 55824 32895
rect 56784 32920 56836 32972
rect 57152 32963 57204 32972
rect 57152 32929 57161 32963
rect 57161 32929 57195 32963
rect 57195 32929 57204 32963
rect 57152 32920 57204 32929
rect 57980 32920 58032 32972
rect 55772 32852 55824 32861
rect 56232 32852 56284 32904
rect 57060 32784 57112 32836
rect 57428 32852 57480 32904
rect 58256 32784 58308 32836
rect 44456 32759 44508 32768
rect 44456 32725 44465 32759
rect 44465 32725 44499 32759
rect 44499 32725 44508 32759
rect 44456 32716 44508 32725
rect 45284 32759 45336 32768
rect 45284 32725 45293 32759
rect 45293 32725 45327 32759
rect 45327 32725 45336 32759
rect 45284 32716 45336 32725
rect 47952 32716 48004 32768
rect 48596 32716 48648 32768
rect 52736 32716 52788 32768
rect 58164 32716 58216 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 29736 32512 29788 32564
rect 30288 32512 30340 32564
rect 28356 32487 28408 32496
rect 28356 32453 28365 32487
rect 28365 32453 28399 32487
rect 28399 32453 28408 32487
rect 28356 32444 28408 32453
rect 29644 32444 29696 32496
rect 30196 32444 30248 32496
rect 31024 32512 31076 32564
rect 31576 32512 31628 32564
rect 32864 32512 32916 32564
rect 34704 32555 34756 32564
rect 34244 32444 34296 32496
rect 34704 32521 34713 32555
rect 34713 32521 34747 32555
rect 34747 32521 34756 32555
rect 34704 32512 34756 32521
rect 35808 32512 35860 32564
rect 36084 32512 36136 32564
rect 32312 32308 32364 32360
rect 34888 32376 34940 32428
rect 35532 32376 35584 32428
rect 32956 32351 33008 32360
rect 32956 32317 32965 32351
rect 32965 32317 32999 32351
rect 32999 32317 33008 32351
rect 32956 32308 33008 32317
rect 37372 32512 37424 32564
rect 37556 32555 37608 32564
rect 37556 32521 37565 32555
rect 37565 32521 37599 32555
rect 37599 32521 37608 32555
rect 37556 32512 37608 32521
rect 38200 32512 38252 32564
rect 38614 32512 38666 32564
rect 39120 32555 39172 32564
rect 37280 32444 37332 32496
rect 37924 32444 37976 32496
rect 38844 32444 38896 32496
rect 39120 32521 39129 32555
rect 39129 32521 39163 32555
rect 39163 32521 39172 32555
rect 39120 32512 39172 32521
rect 40408 32512 40460 32564
rect 36544 32308 36596 32360
rect 36452 32240 36504 32292
rect 36912 32351 36964 32360
rect 36912 32317 36921 32351
rect 36921 32317 36955 32351
rect 36955 32317 36964 32351
rect 36912 32308 36964 32317
rect 38476 32419 38528 32428
rect 38476 32385 38511 32419
rect 38511 32385 38528 32419
rect 38476 32376 38528 32385
rect 38660 32419 38712 32428
rect 38660 32385 38669 32419
rect 38669 32385 38703 32419
rect 38703 32385 38712 32419
rect 39304 32419 39356 32428
rect 38660 32376 38712 32385
rect 39304 32385 39313 32419
rect 39313 32385 39347 32419
rect 39347 32385 39356 32419
rect 39304 32376 39356 32385
rect 39212 32308 39264 32360
rect 39580 32419 39632 32428
rect 41604 32512 41656 32564
rect 42892 32512 42944 32564
rect 43720 32512 43772 32564
rect 46940 32512 46992 32564
rect 47216 32555 47268 32564
rect 47216 32521 47225 32555
rect 47225 32521 47259 32555
rect 47259 32521 47268 32555
rect 47216 32512 47268 32521
rect 49792 32512 49844 32564
rect 50804 32512 50856 32564
rect 39580 32385 39615 32419
rect 39615 32385 39632 32419
rect 39580 32376 39632 32385
rect 40408 32419 40460 32428
rect 40408 32385 40417 32419
rect 40417 32385 40451 32419
rect 40451 32385 40460 32419
rect 40408 32376 40460 32385
rect 40592 32419 40644 32428
rect 40592 32385 40601 32419
rect 40601 32385 40635 32419
rect 40635 32385 40644 32419
rect 40592 32376 40644 32385
rect 41328 32376 41380 32428
rect 35348 32172 35400 32224
rect 36268 32172 36320 32224
rect 37556 32172 37608 32224
rect 39580 32240 39632 32292
rect 39856 32308 39908 32360
rect 41236 32240 41288 32292
rect 39212 32172 39264 32224
rect 40224 32172 40276 32224
rect 44456 32444 44508 32496
rect 42800 32419 42852 32428
rect 42800 32385 42809 32419
rect 42809 32385 42843 32419
rect 42843 32385 42852 32419
rect 42800 32376 42852 32385
rect 42984 32419 43036 32428
rect 42984 32385 42993 32419
rect 42993 32385 43027 32419
rect 43027 32385 43036 32419
rect 42984 32376 43036 32385
rect 43720 32419 43772 32428
rect 43720 32385 43729 32419
rect 43729 32385 43763 32419
rect 43763 32385 43772 32419
rect 43720 32376 43772 32385
rect 45928 32444 45980 32496
rect 48412 32444 48464 32496
rect 46848 32376 46900 32428
rect 48596 32376 48648 32428
rect 49424 32444 49476 32496
rect 51356 32512 51408 32564
rect 52000 32512 52052 32564
rect 52736 32512 52788 32564
rect 52920 32555 52972 32564
rect 52920 32521 52929 32555
rect 52929 32521 52963 32555
rect 52963 32521 52972 32555
rect 52920 32512 52972 32521
rect 53932 32512 53984 32564
rect 56232 32555 56284 32564
rect 56232 32521 56241 32555
rect 56241 32521 56275 32555
rect 56275 32521 56284 32555
rect 56232 32512 56284 32521
rect 57152 32512 57204 32564
rect 50712 32419 50764 32428
rect 50712 32385 50721 32419
rect 50721 32385 50755 32419
rect 50755 32385 50764 32419
rect 50712 32376 50764 32385
rect 46020 32308 46072 32360
rect 47124 32308 47176 32360
rect 50896 32419 50948 32428
rect 50896 32385 50905 32419
rect 50905 32385 50939 32419
rect 50939 32385 50948 32419
rect 50896 32376 50948 32385
rect 51080 32419 51132 32428
rect 51080 32385 51089 32419
rect 51089 32385 51123 32419
rect 51123 32385 51132 32419
rect 51080 32376 51132 32385
rect 51632 32376 51684 32428
rect 51908 32419 51960 32428
rect 51908 32385 51917 32419
rect 51917 32385 51951 32419
rect 51951 32385 51960 32419
rect 51908 32376 51960 32385
rect 52000 32419 52052 32428
rect 52000 32385 52045 32419
rect 52045 32385 52052 32419
rect 52000 32376 52052 32385
rect 52184 32419 52236 32428
rect 52184 32385 52193 32419
rect 52193 32385 52227 32419
rect 52227 32385 52236 32419
rect 52184 32376 52236 32385
rect 52644 32376 52696 32428
rect 53380 32444 53432 32496
rect 54392 32444 54444 32496
rect 54944 32444 54996 32496
rect 55772 32444 55824 32496
rect 50988 32308 51040 32360
rect 52552 32308 52604 32360
rect 53288 32308 53340 32360
rect 52276 32240 52328 32292
rect 53656 32376 53708 32428
rect 54576 32376 54628 32428
rect 55588 32419 55640 32428
rect 55588 32385 55597 32419
rect 55597 32385 55631 32419
rect 55631 32385 55640 32419
rect 55588 32376 55640 32385
rect 54116 32308 54168 32360
rect 55956 32419 56008 32428
rect 55956 32385 55965 32419
rect 55965 32385 55999 32419
rect 55999 32385 56008 32419
rect 55956 32376 56008 32385
rect 56324 32444 56376 32496
rect 56416 32376 56468 32428
rect 56784 32419 56836 32428
rect 56784 32385 56793 32419
rect 56793 32385 56827 32419
rect 56827 32385 56836 32419
rect 57336 32444 57388 32496
rect 56784 32376 56836 32385
rect 57060 32419 57112 32428
rect 57060 32385 57069 32419
rect 57069 32385 57103 32419
rect 57103 32385 57112 32419
rect 57060 32376 57112 32385
rect 55956 32240 56008 32292
rect 48136 32172 48188 32224
rect 49516 32172 49568 32224
rect 52368 32172 52420 32224
rect 52644 32172 52696 32224
rect 53656 32172 53708 32224
rect 57980 32172 58032 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 30288 31968 30340 32020
rect 31116 31968 31168 32020
rect 32312 31968 32364 32020
rect 30196 31900 30248 31952
rect 34244 31968 34296 32020
rect 35348 32011 35400 32020
rect 35348 31977 35357 32011
rect 35357 31977 35391 32011
rect 35391 31977 35400 32011
rect 35348 31968 35400 31977
rect 36360 31968 36412 32020
rect 37280 31968 37332 32020
rect 38476 31968 38528 32020
rect 38568 31968 38620 32020
rect 38660 31968 38712 32020
rect 41236 31968 41288 32020
rect 41604 32011 41656 32020
rect 41604 31977 41613 32011
rect 41613 31977 41647 32011
rect 41647 31977 41656 32011
rect 41604 31968 41656 31977
rect 42892 31968 42944 32020
rect 43904 31968 43956 32020
rect 46940 32011 46992 32020
rect 46940 31977 46949 32011
rect 46949 31977 46983 32011
rect 46983 31977 46992 32011
rect 46940 31968 46992 31977
rect 47768 31968 47820 32020
rect 48136 32011 48188 32020
rect 48136 31977 48145 32011
rect 48145 31977 48179 32011
rect 48179 31977 48188 32011
rect 48136 31968 48188 31977
rect 48688 31968 48740 32020
rect 49056 31968 49108 32020
rect 52184 31968 52236 32020
rect 42432 31900 42484 31952
rect 47584 31900 47636 31952
rect 32956 31875 33008 31884
rect 32956 31841 32965 31875
rect 32965 31841 32999 31875
rect 32999 31841 33008 31875
rect 32956 31832 33008 31841
rect 34612 31832 34664 31884
rect 35348 31832 35400 31884
rect 35532 31832 35584 31884
rect 35900 31832 35952 31884
rect 36084 31832 36136 31884
rect 36268 31832 36320 31884
rect 30288 31764 30340 31816
rect 34704 31764 34756 31816
rect 32404 31696 32456 31748
rect 32680 31739 32732 31748
rect 32680 31705 32689 31739
rect 32689 31705 32723 31739
rect 32723 31705 32732 31739
rect 32680 31696 32732 31705
rect 36544 31764 36596 31816
rect 36728 31807 36780 31816
rect 36728 31773 36737 31807
rect 36737 31773 36771 31807
rect 36771 31773 36780 31807
rect 36728 31764 36780 31773
rect 37280 31832 37332 31884
rect 37188 31807 37240 31816
rect 37188 31773 37197 31807
rect 37197 31773 37231 31807
rect 37231 31773 37240 31807
rect 37188 31764 37240 31773
rect 38292 31832 38344 31884
rect 42156 31875 42208 31884
rect 37556 31764 37608 31816
rect 40224 31807 40276 31816
rect 40224 31773 40233 31807
rect 40233 31773 40267 31807
rect 40267 31773 40276 31807
rect 40224 31764 40276 31773
rect 40408 31807 40460 31816
rect 40408 31773 40417 31807
rect 40417 31773 40451 31807
rect 40451 31773 40460 31807
rect 40408 31764 40460 31773
rect 29828 31671 29880 31680
rect 29828 31637 29837 31671
rect 29837 31637 29871 31671
rect 29871 31637 29880 31671
rect 29828 31628 29880 31637
rect 35808 31628 35860 31680
rect 36268 31628 36320 31680
rect 36820 31628 36872 31680
rect 38844 31696 38896 31748
rect 40040 31696 40092 31748
rect 42156 31841 42165 31875
rect 42165 31841 42199 31875
rect 42199 31841 42208 31875
rect 42156 31832 42208 31841
rect 42892 31832 42944 31884
rect 43260 31832 43312 31884
rect 47216 31832 47268 31884
rect 47676 31832 47728 31884
rect 41328 31764 41380 31816
rect 42800 31764 42852 31816
rect 43076 31764 43128 31816
rect 44272 31807 44324 31816
rect 44272 31773 44281 31807
rect 44281 31773 44315 31807
rect 44315 31773 44324 31807
rect 44272 31764 44324 31773
rect 45928 31807 45980 31816
rect 45928 31773 45937 31807
rect 45937 31773 45971 31807
rect 45971 31773 45980 31807
rect 45928 31764 45980 31773
rect 48228 31807 48280 31816
rect 48228 31773 48237 31807
rect 48237 31773 48271 31807
rect 48271 31773 48280 31807
rect 48228 31764 48280 31773
rect 48596 31764 48648 31816
rect 51908 31900 51960 31952
rect 53380 31968 53432 32020
rect 54484 31968 54536 32020
rect 56416 32011 56468 32020
rect 56416 31977 56425 32011
rect 56425 31977 56459 32011
rect 56459 31977 56468 32011
rect 56416 31968 56468 31977
rect 50896 31832 50948 31884
rect 42892 31696 42944 31748
rect 38936 31628 38988 31680
rect 39028 31628 39080 31680
rect 43076 31671 43128 31680
rect 43076 31637 43085 31671
rect 43085 31637 43119 31671
rect 43119 31637 43128 31671
rect 43076 31628 43128 31637
rect 45560 31696 45612 31748
rect 46020 31739 46072 31748
rect 46020 31705 46029 31739
rect 46029 31705 46063 31739
rect 46063 31705 46072 31739
rect 46020 31696 46072 31705
rect 45284 31628 45336 31680
rect 47860 31696 47912 31748
rect 50988 31807 51040 31816
rect 50988 31773 50997 31807
rect 50997 31773 51031 31807
rect 51031 31773 51040 31807
rect 50988 31764 51040 31773
rect 51448 31807 51500 31816
rect 51448 31773 51457 31807
rect 51457 31773 51491 31807
rect 51491 31773 51500 31807
rect 51448 31764 51500 31773
rect 51632 31807 51684 31816
rect 51632 31773 51641 31807
rect 51641 31773 51675 31807
rect 51675 31773 51684 31807
rect 51632 31764 51684 31773
rect 52552 31807 52604 31816
rect 50804 31739 50856 31748
rect 50804 31705 50813 31739
rect 50813 31705 50847 31739
rect 50847 31705 50856 31739
rect 50804 31696 50856 31705
rect 52552 31773 52561 31807
rect 52561 31773 52595 31807
rect 52595 31773 52604 31807
rect 52552 31764 52604 31773
rect 54576 31900 54628 31952
rect 53288 31807 53340 31816
rect 53288 31773 53295 31807
rect 53295 31773 53340 31807
rect 52368 31696 52420 31748
rect 53288 31764 53340 31773
rect 53564 31807 53616 31816
rect 53564 31773 53578 31807
rect 53578 31773 53612 31807
rect 53612 31773 53616 31807
rect 53564 31764 53616 31773
rect 54944 31764 54996 31816
rect 55404 31832 55456 31884
rect 55588 31764 55640 31816
rect 54392 31696 54444 31748
rect 56324 31832 56376 31884
rect 55956 31764 56008 31816
rect 56140 31807 56192 31816
rect 56140 31773 56149 31807
rect 56149 31773 56183 31807
rect 56183 31773 56192 31807
rect 56140 31764 56192 31773
rect 58072 31900 58124 31952
rect 58348 31832 58400 31884
rect 57612 31807 57664 31816
rect 57612 31773 57621 31807
rect 57621 31773 57655 31807
rect 57655 31773 57664 31807
rect 57612 31764 57664 31773
rect 58256 31764 58308 31816
rect 58532 31764 58584 31816
rect 57796 31696 57848 31748
rect 46388 31671 46440 31680
rect 46388 31637 46397 31671
rect 46397 31637 46431 31671
rect 46431 31637 46440 31671
rect 46388 31628 46440 31637
rect 47124 31628 47176 31680
rect 47584 31628 47636 31680
rect 55036 31628 55088 31680
rect 57980 31628 58032 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 28264 31424 28316 31476
rect 32404 31467 32456 31476
rect 32404 31433 32413 31467
rect 32413 31433 32447 31467
rect 32447 31433 32456 31467
rect 32404 31424 32456 31433
rect 32680 31424 32732 31476
rect 29828 31356 29880 31408
rect 33876 31356 33928 31408
rect 34612 31356 34664 31408
rect 30196 31331 30248 31340
rect 30196 31297 30205 31331
rect 30205 31297 30239 31331
rect 30239 31297 30248 31331
rect 30196 31288 30248 31297
rect 32864 31288 32916 31340
rect 32956 31288 33008 31340
rect 35348 31424 35400 31476
rect 36268 31424 36320 31476
rect 38108 31467 38160 31476
rect 38108 31433 38117 31467
rect 38117 31433 38151 31467
rect 38151 31433 38160 31467
rect 38108 31424 38160 31433
rect 39856 31424 39908 31476
rect 38844 31399 38896 31408
rect 38844 31365 38871 31399
rect 38871 31365 38896 31399
rect 38844 31356 38896 31365
rect 39028 31399 39080 31408
rect 39028 31365 39037 31399
rect 39037 31365 39071 31399
rect 39071 31365 39080 31399
rect 39028 31356 39080 31365
rect 33692 31220 33744 31272
rect 33968 31084 34020 31136
rect 35808 31084 35860 31136
rect 36084 31263 36136 31272
rect 36084 31229 36093 31263
rect 36093 31229 36127 31263
rect 36127 31229 36136 31263
rect 36452 31288 36504 31340
rect 39488 31356 39540 31408
rect 40316 31424 40368 31476
rect 41328 31424 41380 31476
rect 45928 31424 45980 31476
rect 40592 31356 40644 31408
rect 46020 31399 46072 31408
rect 46020 31365 46029 31399
rect 46029 31365 46063 31399
rect 46063 31365 46072 31399
rect 46020 31356 46072 31365
rect 39304 31288 39356 31340
rect 39764 31288 39816 31340
rect 36084 31220 36136 31229
rect 40040 31220 40092 31272
rect 40868 31288 40920 31340
rect 41512 31331 41564 31340
rect 41512 31297 41521 31331
rect 41521 31297 41555 31331
rect 41555 31297 41564 31331
rect 41512 31288 41564 31297
rect 43352 31331 43404 31340
rect 43352 31297 43361 31331
rect 43361 31297 43395 31331
rect 43395 31297 43404 31331
rect 43352 31288 43404 31297
rect 43720 31288 43772 31340
rect 44088 31331 44140 31340
rect 44088 31297 44097 31331
rect 44097 31297 44131 31331
rect 44131 31297 44140 31331
rect 44088 31288 44140 31297
rect 45192 31331 45244 31340
rect 45192 31297 45201 31331
rect 45201 31297 45235 31331
rect 45235 31297 45244 31331
rect 48320 31424 48372 31476
rect 46848 31356 46900 31408
rect 47676 31356 47728 31408
rect 50988 31424 51040 31476
rect 52644 31424 52696 31476
rect 46940 31331 46992 31340
rect 45192 31288 45244 31297
rect 46940 31297 46949 31331
rect 46949 31297 46983 31331
rect 46983 31297 46992 31331
rect 46940 31288 46992 31297
rect 37004 31152 37056 31204
rect 39028 31152 39080 31204
rect 42892 31220 42944 31272
rect 42984 31220 43036 31272
rect 44640 31220 44692 31272
rect 46204 31220 46256 31272
rect 48320 31288 48372 31340
rect 50804 31331 50856 31340
rect 48964 31263 49016 31272
rect 42432 31152 42484 31204
rect 42708 31195 42760 31204
rect 42708 31161 42717 31195
rect 42717 31161 42751 31195
rect 42751 31161 42760 31195
rect 42708 31152 42760 31161
rect 43168 31195 43220 31204
rect 43168 31161 43177 31195
rect 43177 31161 43211 31195
rect 43211 31161 43220 31195
rect 43168 31152 43220 31161
rect 47216 31152 47268 31204
rect 37464 31084 37516 31136
rect 38752 31084 38804 31136
rect 41788 31084 41840 31136
rect 43444 31084 43496 31136
rect 46940 31127 46992 31136
rect 46940 31093 46949 31127
rect 46949 31093 46983 31127
rect 46983 31093 46992 31127
rect 46940 31084 46992 31093
rect 47032 31084 47084 31136
rect 48964 31229 48973 31263
rect 48973 31229 49007 31263
rect 49007 31229 49016 31263
rect 48964 31220 49016 31229
rect 48412 31152 48464 31204
rect 50804 31297 50814 31331
rect 50814 31297 50856 31331
rect 50804 31288 50856 31297
rect 51908 31356 51960 31408
rect 51540 31331 51592 31340
rect 51540 31297 51549 31331
rect 51549 31297 51583 31331
rect 51583 31297 51592 31331
rect 51540 31288 51592 31297
rect 53564 31356 53616 31408
rect 54116 31356 54168 31408
rect 53748 31288 53800 31340
rect 54300 31288 54352 31340
rect 54484 31331 54536 31340
rect 54484 31297 54493 31331
rect 54493 31297 54527 31331
rect 54527 31297 54536 31331
rect 54484 31288 54536 31297
rect 54576 31331 54628 31340
rect 54576 31297 54585 31331
rect 54585 31297 54619 31331
rect 54619 31297 54628 31331
rect 54576 31288 54628 31297
rect 55036 31288 55088 31340
rect 56324 31356 56376 31408
rect 56140 31331 56192 31340
rect 50344 31195 50396 31204
rect 50344 31161 50353 31195
rect 50353 31161 50387 31195
rect 50387 31161 50396 31195
rect 50344 31152 50396 31161
rect 49608 31084 49660 31136
rect 49884 31084 49936 31136
rect 54116 31263 54168 31272
rect 54116 31229 54125 31263
rect 54125 31229 54159 31263
rect 54159 31229 54168 31263
rect 54116 31220 54168 31229
rect 54392 31220 54444 31272
rect 55588 31220 55640 31272
rect 56140 31297 56149 31331
rect 56149 31297 56183 31331
rect 56183 31297 56192 31331
rect 56140 31288 56192 31297
rect 56784 31356 56836 31408
rect 57060 31356 57112 31408
rect 58532 31288 58584 31340
rect 57888 31220 57940 31272
rect 58072 31263 58124 31272
rect 58072 31229 58081 31263
rect 58081 31229 58115 31263
rect 58115 31229 58124 31263
rect 58072 31220 58124 31229
rect 57612 31152 57664 31204
rect 51356 31127 51408 31136
rect 51356 31093 51365 31127
rect 51365 31093 51399 31127
rect 51399 31093 51408 31127
rect 51356 31084 51408 31093
rect 52276 31084 52328 31136
rect 53380 31084 53432 31136
rect 54760 31127 54812 31136
rect 54760 31093 54769 31127
rect 54769 31093 54803 31127
rect 54803 31093 54812 31127
rect 54760 31084 54812 31093
rect 57152 31084 57204 31136
rect 57796 31084 57848 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 33692 30923 33744 30932
rect 33692 30889 33701 30923
rect 33701 30889 33735 30923
rect 33735 30889 33744 30923
rect 33692 30880 33744 30889
rect 38752 30880 38804 30932
rect 40408 30880 40460 30932
rect 44272 30880 44324 30932
rect 46572 30880 46624 30932
rect 33876 30812 33928 30864
rect 29460 30744 29512 30796
rect 34796 30744 34848 30796
rect 35348 30744 35400 30796
rect 39396 30812 39448 30864
rect 51540 30880 51592 30932
rect 43352 30744 43404 30796
rect 31852 30719 31904 30728
rect 31852 30685 31861 30719
rect 31861 30685 31895 30719
rect 31895 30685 31904 30719
rect 31852 30676 31904 30685
rect 30840 30608 30892 30660
rect 31668 30608 31720 30660
rect 33968 30676 34020 30728
rect 34152 30676 34204 30728
rect 39764 30676 39816 30728
rect 40408 30719 40460 30728
rect 40408 30685 40417 30719
rect 40417 30685 40451 30719
rect 40451 30685 40460 30719
rect 40408 30676 40460 30685
rect 40776 30676 40828 30728
rect 41328 30676 41380 30728
rect 43076 30676 43128 30728
rect 43904 30676 43956 30728
rect 1676 30583 1728 30592
rect 1676 30549 1685 30583
rect 1685 30549 1719 30583
rect 1719 30549 1728 30583
rect 1676 30540 1728 30549
rect 2412 30583 2464 30592
rect 2412 30549 2421 30583
rect 2421 30549 2455 30583
rect 2455 30549 2464 30583
rect 2412 30540 2464 30549
rect 34796 30540 34848 30592
rect 36176 30608 36228 30660
rect 36360 30608 36412 30660
rect 35164 30540 35216 30592
rect 35808 30540 35860 30592
rect 36452 30540 36504 30592
rect 37464 30608 37516 30660
rect 38936 30651 38988 30660
rect 38936 30617 38945 30651
rect 38945 30617 38979 30651
rect 38979 30617 38988 30651
rect 38936 30608 38988 30617
rect 40040 30608 40092 30660
rect 40316 30651 40368 30660
rect 40316 30617 40325 30651
rect 40325 30617 40359 30651
rect 40359 30617 40368 30651
rect 40316 30608 40368 30617
rect 40500 30651 40552 30660
rect 40500 30617 40535 30651
rect 40535 30617 40552 30651
rect 41788 30651 41840 30660
rect 40500 30608 40552 30617
rect 41788 30617 41797 30651
rect 41797 30617 41831 30651
rect 41831 30617 41840 30651
rect 41788 30608 41840 30617
rect 43444 30608 43496 30660
rect 43720 30608 43772 30660
rect 45284 30608 45336 30660
rect 45928 30676 45980 30728
rect 46112 30676 46164 30728
rect 46572 30676 46624 30728
rect 46756 30719 46808 30728
rect 46756 30685 46765 30719
rect 46765 30685 46799 30719
rect 46799 30685 46808 30719
rect 47584 30719 47636 30728
rect 46756 30676 46808 30685
rect 47584 30685 47593 30719
rect 47593 30685 47627 30719
rect 47627 30685 47636 30719
rect 47584 30676 47636 30685
rect 48412 30744 48464 30796
rect 50988 30812 51040 30864
rect 55864 30880 55916 30932
rect 57612 30880 57664 30932
rect 54024 30812 54076 30864
rect 50344 30744 50396 30796
rect 50804 30744 50856 30796
rect 47860 30719 47912 30728
rect 47860 30685 47895 30719
rect 47895 30685 47912 30719
rect 48044 30719 48096 30728
rect 47860 30676 47912 30685
rect 48044 30685 48053 30719
rect 48053 30685 48087 30719
rect 48087 30685 48096 30719
rect 48044 30676 48096 30685
rect 49056 30719 49108 30728
rect 49056 30685 49065 30719
rect 49065 30685 49099 30719
rect 49099 30685 49108 30719
rect 49056 30676 49108 30685
rect 51448 30744 51500 30796
rect 52460 30787 52512 30796
rect 52460 30753 52469 30787
rect 52469 30753 52503 30787
rect 52503 30753 52512 30787
rect 52460 30744 52512 30753
rect 52736 30744 52788 30796
rect 54300 30812 54352 30864
rect 54576 30812 54628 30864
rect 51172 30719 51224 30728
rect 38844 30540 38896 30592
rect 44180 30583 44232 30592
rect 44180 30549 44189 30583
rect 44189 30549 44223 30583
rect 44223 30549 44232 30583
rect 44180 30540 44232 30549
rect 46020 30540 46072 30592
rect 46848 30540 46900 30592
rect 47584 30540 47636 30592
rect 47676 30540 47728 30592
rect 48136 30608 48188 30660
rect 49700 30608 49752 30660
rect 50620 30608 50672 30660
rect 51172 30685 51181 30719
rect 51181 30685 51215 30719
rect 51215 30685 51224 30719
rect 51172 30676 51224 30685
rect 51632 30676 51684 30728
rect 52552 30719 52604 30728
rect 52552 30685 52561 30719
rect 52561 30685 52595 30719
rect 52595 30685 52604 30719
rect 52552 30676 52604 30685
rect 54484 30676 54536 30728
rect 54760 30676 54812 30728
rect 57336 30744 57388 30796
rect 58440 30744 58492 30796
rect 57152 30719 57204 30728
rect 52000 30608 52052 30660
rect 52184 30608 52236 30660
rect 52828 30651 52880 30660
rect 52368 30540 52420 30592
rect 52828 30617 52837 30651
rect 52837 30617 52871 30651
rect 52871 30617 52880 30651
rect 52828 30608 52880 30617
rect 54116 30608 54168 30660
rect 54576 30651 54628 30660
rect 54576 30617 54585 30651
rect 54585 30617 54619 30651
rect 54619 30617 54628 30651
rect 54576 30608 54628 30617
rect 53840 30540 53892 30592
rect 54944 30608 54996 30660
rect 57152 30685 57161 30719
rect 57161 30685 57195 30719
rect 57195 30685 57204 30719
rect 57152 30676 57204 30685
rect 56508 30608 56560 30660
rect 57060 30540 57112 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 34704 30336 34756 30388
rect 34796 30336 34848 30388
rect 30840 30311 30892 30320
rect 30840 30277 30849 30311
rect 30849 30277 30883 30311
rect 30883 30277 30892 30311
rect 30840 30268 30892 30277
rect 35164 30336 35216 30388
rect 35624 30336 35676 30388
rect 36360 30379 36412 30388
rect 36360 30345 36369 30379
rect 36369 30345 36403 30379
rect 36403 30345 36412 30379
rect 36360 30336 36412 30345
rect 36728 30336 36780 30388
rect 37280 30336 37332 30388
rect 35348 30268 35400 30320
rect 37556 30268 37608 30320
rect 37924 30311 37976 30320
rect 37924 30277 37959 30311
rect 37959 30277 37976 30311
rect 37924 30268 37976 30277
rect 38568 30268 38620 30320
rect 28816 30243 28868 30252
rect 28816 30209 28825 30243
rect 28825 30209 28859 30243
rect 28859 30209 28868 30243
rect 28816 30200 28868 30209
rect 28908 30200 28960 30252
rect 30288 30200 30340 30252
rect 31760 30200 31812 30252
rect 32772 30200 32824 30252
rect 34152 30243 34204 30252
rect 34152 30209 34161 30243
rect 34161 30209 34195 30243
rect 34195 30209 34204 30243
rect 34152 30200 34204 30209
rect 40040 30311 40092 30320
rect 40040 30277 40049 30311
rect 40049 30277 40083 30311
rect 40083 30277 40092 30311
rect 41052 30336 41104 30388
rect 40040 30268 40092 30277
rect 37832 30243 37884 30252
rect 37832 30209 37842 30243
rect 37842 30209 37876 30243
rect 37876 30209 37884 30243
rect 37832 30200 37884 30209
rect 28540 30064 28592 30116
rect 31760 29996 31812 30048
rect 32404 30039 32456 30048
rect 32404 30005 32413 30039
rect 32413 30005 32447 30039
rect 32447 30005 32456 30039
rect 32404 29996 32456 30005
rect 34888 30132 34940 30184
rect 38108 30243 38160 30252
rect 38108 30209 38117 30243
rect 38117 30209 38151 30243
rect 38151 30209 38160 30243
rect 38108 30200 38160 30209
rect 38660 30200 38712 30252
rect 39948 30243 40000 30252
rect 39028 30132 39080 30184
rect 39948 30209 39957 30243
rect 39957 30209 39991 30243
rect 39991 30209 40000 30243
rect 39948 30200 40000 30209
rect 39212 30132 39264 30184
rect 40684 30268 40736 30320
rect 40868 30268 40920 30320
rect 45192 30311 45244 30320
rect 45192 30277 45201 30311
rect 45201 30277 45235 30311
rect 45235 30277 45244 30311
rect 45192 30268 45244 30277
rect 45744 30268 45796 30320
rect 47676 30336 47728 30388
rect 48320 30336 48372 30388
rect 40500 30200 40552 30252
rect 41512 30243 41564 30252
rect 41512 30209 41520 30243
rect 41520 30209 41554 30243
rect 41554 30209 41564 30243
rect 41512 30200 41564 30209
rect 42800 30200 42852 30252
rect 43168 30243 43220 30252
rect 43168 30209 43177 30243
rect 43177 30209 43211 30243
rect 43211 30209 43220 30243
rect 43168 30200 43220 30209
rect 44548 30200 44600 30252
rect 45560 30200 45612 30252
rect 49700 30311 49752 30320
rect 49700 30277 49709 30311
rect 49709 30277 49743 30311
rect 49743 30277 49752 30311
rect 49700 30268 49752 30277
rect 50436 30268 50488 30320
rect 46664 30243 46716 30252
rect 46664 30209 46673 30243
rect 46673 30209 46707 30243
rect 46707 30209 46716 30243
rect 46664 30200 46716 30209
rect 46848 30200 46900 30252
rect 40408 30175 40460 30184
rect 35900 30064 35952 30116
rect 40408 30141 40417 30175
rect 40417 30141 40451 30175
rect 40451 30141 40460 30175
rect 40408 30132 40460 30141
rect 40316 30064 40368 30116
rect 40684 30064 40736 30116
rect 40868 30064 40920 30116
rect 41328 30132 41380 30184
rect 45284 30132 45336 30184
rect 47676 30132 47728 30184
rect 48320 30200 48372 30252
rect 42984 30064 43036 30116
rect 46296 30064 46348 30116
rect 48872 30200 48924 30252
rect 51172 30336 51224 30388
rect 52184 30336 52236 30388
rect 50620 30311 50672 30320
rect 50620 30277 50629 30311
rect 50629 30277 50663 30311
rect 50663 30277 50672 30311
rect 50620 30268 50672 30277
rect 48504 30132 48556 30184
rect 50804 30243 50856 30252
rect 50804 30209 50813 30243
rect 50813 30209 50847 30243
rect 50847 30209 50856 30243
rect 50804 30200 50856 30209
rect 52000 30243 52052 30252
rect 52000 30209 52009 30243
rect 52009 30209 52043 30243
rect 52043 30209 52052 30243
rect 52000 30200 52052 30209
rect 52184 30200 52236 30252
rect 53380 30336 53432 30388
rect 52368 30243 52420 30252
rect 52368 30209 52377 30243
rect 52377 30209 52411 30243
rect 52411 30209 52420 30243
rect 52368 30200 52420 30209
rect 53840 30268 53892 30320
rect 49148 30175 49200 30184
rect 49148 30141 49157 30175
rect 49157 30141 49191 30175
rect 49191 30141 49200 30175
rect 53748 30243 53800 30252
rect 53748 30209 53757 30243
rect 53757 30209 53791 30243
rect 53791 30209 53800 30243
rect 53932 30243 53984 30252
rect 53748 30200 53800 30209
rect 53932 30209 53941 30243
rect 53941 30209 53975 30243
rect 53975 30209 53984 30243
rect 53932 30200 53984 30209
rect 54116 30336 54168 30388
rect 57888 30336 57940 30388
rect 55036 30268 55088 30320
rect 55312 30268 55364 30320
rect 56600 30268 56652 30320
rect 54208 30200 54260 30252
rect 54944 30200 54996 30252
rect 55772 30200 55824 30252
rect 56140 30200 56192 30252
rect 57336 30200 57388 30252
rect 49148 30132 49200 30141
rect 53288 30132 53340 30184
rect 55496 30132 55548 30184
rect 56416 30175 56468 30184
rect 52552 30064 52604 30116
rect 56416 30141 56425 30175
rect 56425 30141 56459 30175
rect 56459 30141 56468 30175
rect 56416 30132 56468 30141
rect 57060 30175 57112 30184
rect 57060 30141 57069 30175
rect 57069 30141 57103 30175
rect 57103 30141 57112 30175
rect 57060 30132 57112 30141
rect 56048 30064 56100 30116
rect 57520 30107 57572 30116
rect 57520 30073 57529 30107
rect 57529 30073 57563 30107
rect 57563 30073 57572 30107
rect 57520 30064 57572 30073
rect 34520 29996 34572 30048
rect 34704 29996 34756 30048
rect 35440 29996 35492 30048
rect 35532 29996 35584 30048
rect 38200 29996 38252 30048
rect 38476 29996 38528 30048
rect 41512 29996 41564 30048
rect 41604 29996 41656 30048
rect 50252 29996 50304 30048
rect 51908 29996 51960 30048
rect 53104 29996 53156 30048
rect 53564 29996 53616 30048
rect 55128 29996 55180 30048
rect 55956 29996 56008 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 29368 29792 29420 29844
rect 31852 29792 31904 29844
rect 33416 29792 33468 29844
rect 34152 29792 34204 29844
rect 35348 29792 35400 29844
rect 36452 29835 36504 29844
rect 36452 29801 36461 29835
rect 36461 29801 36495 29835
rect 36495 29801 36504 29835
rect 36452 29792 36504 29801
rect 30196 29588 30248 29640
rect 31668 29588 31720 29640
rect 35900 29724 35952 29776
rect 37556 29767 37608 29776
rect 31300 29563 31352 29572
rect 31300 29529 31309 29563
rect 31309 29529 31343 29563
rect 31343 29529 31352 29563
rect 31300 29520 31352 29529
rect 32956 29520 33008 29572
rect 28816 29452 28868 29504
rect 34796 29588 34848 29640
rect 35532 29588 35584 29640
rect 37556 29733 37565 29767
rect 37565 29733 37599 29767
rect 37599 29733 37608 29767
rect 37556 29724 37608 29733
rect 38568 29724 38620 29776
rect 39764 29724 39816 29776
rect 40132 29724 40184 29776
rect 40408 29724 40460 29776
rect 37372 29656 37424 29708
rect 38936 29656 38988 29708
rect 41788 29792 41840 29844
rect 42708 29792 42760 29844
rect 44548 29835 44600 29844
rect 44548 29801 44557 29835
rect 44557 29801 44591 29835
rect 44591 29801 44600 29835
rect 44548 29792 44600 29801
rect 46388 29835 46440 29844
rect 46388 29801 46397 29835
rect 46397 29801 46431 29835
rect 46431 29801 46440 29835
rect 46388 29792 46440 29801
rect 46664 29792 46716 29844
rect 47216 29835 47268 29844
rect 47216 29801 47225 29835
rect 47225 29801 47259 29835
rect 47259 29801 47268 29835
rect 47216 29792 47268 29801
rect 47676 29792 47728 29844
rect 49148 29792 49200 29844
rect 53748 29792 53800 29844
rect 41328 29724 41380 29776
rect 47584 29724 47636 29776
rect 49056 29724 49108 29776
rect 42800 29656 42852 29708
rect 44272 29656 44324 29708
rect 36820 29631 36872 29640
rect 36820 29597 36829 29631
rect 36829 29597 36863 29631
rect 36863 29597 36872 29631
rect 36820 29588 36872 29597
rect 34336 29563 34388 29572
rect 34336 29529 34345 29563
rect 34345 29529 34379 29563
rect 34379 29529 34388 29563
rect 34336 29520 34388 29529
rect 35992 29520 36044 29572
rect 34612 29452 34664 29504
rect 35164 29452 35216 29504
rect 35256 29452 35308 29504
rect 35624 29452 35676 29504
rect 36912 29563 36964 29572
rect 36912 29529 36947 29563
rect 36947 29529 36964 29563
rect 36912 29520 36964 29529
rect 37280 29452 37332 29504
rect 38660 29588 38712 29640
rect 40132 29588 40184 29640
rect 41880 29588 41932 29640
rect 43352 29588 43404 29640
rect 43996 29631 44048 29640
rect 43996 29597 44005 29631
rect 44005 29597 44039 29631
rect 44039 29597 44048 29631
rect 43996 29588 44048 29597
rect 44088 29588 44140 29640
rect 45192 29631 45244 29640
rect 45192 29597 45201 29631
rect 45201 29597 45235 29631
rect 45235 29597 45244 29631
rect 45192 29588 45244 29597
rect 45284 29631 45336 29640
rect 45284 29597 45294 29631
rect 45294 29597 45328 29631
rect 45328 29597 45336 29631
rect 46112 29656 46164 29708
rect 46848 29656 46900 29708
rect 47032 29699 47084 29708
rect 47032 29665 47041 29699
rect 47041 29665 47075 29699
rect 47075 29665 47084 29699
rect 47032 29656 47084 29665
rect 47216 29656 47268 29708
rect 51908 29699 51960 29708
rect 51908 29665 51917 29699
rect 51917 29665 51951 29699
rect 51951 29665 51960 29699
rect 51908 29656 51960 29665
rect 53564 29656 53616 29708
rect 56508 29724 56560 29776
rect 56876 29724 56928 29776
rect 54668 29656 54720 29708
rect 55128 29656 55180 29708
rect 45284 29588 45336 29597
rect 46664 29588 46716 29640
rect 47400 29588 47452 29640
rect 47952 29588 48004 29640
rect 41604 29520 41656 29572
rect 41696 29520 41748 29572
rect 43812 29520 43864 29572
rect 45468 29563 45520 29572
rect 45468 29529 45477 29563
rect 45477 29529 45511 29563
rect 45511 29529 45520 29563
rect 45468 29520 45520 29529
rect 45744 29520 45796 29572
rect 47860 29563 47912 29572
rect 47860 29529 47869 29563
rect 47869 29529 47903 29563
rect 47903 29529 47912 29563
rect 47860 29520 47912 29529
rect 48136 29631 48188 29640
rect 48136 29597 48145 29631
rect 48145 29597 48179 29631
rect 48179 29597 48188 29631
rect 48136 29588 48188 29597
rect 48504 29588 48556 29640
rect 48320 29520 48372 29572
rect 50160 29588 50212 29640
rect 38936 29452 38988 29504
rect 40500 29452 40552 29504
rect 42524 29452 42576 29504
rect 43076 29452 43128 29504
rect 48688 29452 48740 29504
rect 49424 29520 49476 29572
rect 52092 29588 52144 29640
rect 52828 29588 52880 29640
rect 53104 29631 53156 29640
rect 53104 29597 53113 29631
rect 53113 29597 53147 29631
rect 53147 29597 53156 29631
rect 53104 29588 53156 29597
rect 53380 29631 53432 29640
rect 53380 29597 53389 29631
rect 53389 29597 53423 29631
rect 53423 29597 53432 29631
rect 53380 29588 53432 29597
rect 53564 29520 53616 29572
rect 49700 29452 49752 29504
rect 49792 29452 49844 29504
rect 52828 29452 52880 29504
rect 53288 29452 53340 29504
rect 55496 29588 55548 29640
rect 55588 29588 55640 29640
rect 55772 29631 55824 29640
rect 55772 29597 55781 29631
rect 55781 29597 55815 29631
rect 55815 29597 55824 29631
rect 56048 29631 56100 29640
rect 55772 29588 55824 29597
rect 56048 29597 56057 29631
rect 56057 29597 56091 29631
rect 56091 29597 56100 29631
rect 56048 29588 56100 29597
rect 57244 29699 57296 29708
rect 57244 29665 57253 29699
rect 57253 29665 57287 29699
rect 57287 29665 57296 29699
rect 57244 29656 57296 29665
rect 57980 29588 58032 29640
rect 55312 29520 55364 29572
rect 56416 29520 56468 29572
rect 55496 29495 55548 29504
rect 55496 29461 55505 29495
rect 55505 29461 55539 29495
rect 55539 29461 55548 29495
rect 55496 29452 55548 29461
rect 58256 29495 58308 29504
rect 58256 29461 58265 29495
rect 58265 29461 58299 29495
rect 58299 29461 58308 29495
rect 58256 29452 58308 29461
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 30196 29291 30248 29300
rect 30196 29257 30205 29291
rect 30205 29257 30239 29291
rect 30239 29257 30248 29291
rect 30196 29248 30248 29257
rect 32772 29248 32824 29300
rect 31760 29155 31812 29164
rect 31760 29121 31769 29155
rect 31769 29121 31803 29155
rect 31803 29121 31812 29155
rect 31760 29112 31812 29121
rect 32864 29112 32916 29164
rect 33416 29155 33468 29164
rect 33416 29121 33425 29155
rect 33425 29121 33459 29155
rect 33459 29121 33468 29155
rect 33416 29112 33468 29121
rect 34796 29112 34848 29164
rect 36820 29248 36872 29300
rect 37372 29248 37424 29300
rect 37648 29248 37700 29300
rect 39212 29291 39264 29300
rect 39212 29257 39221 29291
rect 39221 29257 39255 29291
rect 39255 29257 39264 29291
rect 39212 29248 39264 29257
rect 36360 29180 36412 29232
rect 40040 29248 40092 29300
rect 41144 29248 41196 29300
rect 41696 29291 41748 29300
rect 40776 29180 40828 29232
rect 40868 29180 40920 29232
rect 41420 29223 41472 29232
rect 41420 29189 41429 29223
rect 41429 29189 41463 29223
rect 41463 29189 41472 29223
rect 41420 29180 41472 29189
rect 33692 29087 33744 29096
rect 33692 29053 33701 29087
rect 33701 29053 33735 29087
rect 33735 29053 33744 29087
rect 33692 29044 33744 29053
rect 33784 29044 33836 29096
rect 36912 29112 36964 29164
rect 37556 29112 37608 29164
rect 38844 29155 38896 29164
rect 38844 29121 38853 29155
rect 38853 29121 38887 29155
rect 38887 29121 38896 29155
rect 38844 29112 38896 29121
rect 36360 29087 36412 29096
rect 36360 29053 36369 29087
rect 36369 29053 36403 29087
rect 36403 29053 36412 29087
rect 36360 29044 36412 29053
rect 38568 29044 38620 29096
rect 38936 29044 38988 29096
rect 39948 29112 40000 29164
rect 40316 29112 40368 29164
rect 40500 29155 40552 29164
rect 40500 29121 40509 29155
rect 40509 29121 40543 29155
rect 40543 29121 40552 29155
rect 41052 29155 41104 29164
rect 40500 29112 40552 29121
rect 41052 29121 41061 29155
rect 41061 29121 41095 29155
rect 41095 29121 41104 29155
rect 41052 29112 41104 29121
rect 41236 29155 41288 29164
rect 41236 29121 41253 29155
rect 41253 29121 41288 29155
rect 41236 29112 41288 29121
rect 41696 29257 41705 29291
rect 41705 29257 41739 29291
rect 41739 29257 41748 29291
rect 41696 29248 41748 29257
rect 43352 29248 43404 29300
rect 41880 29180 41932 29232
rect 35164 29019 35216 29028
rect 35164 28985 35173 29019
rect 35173 28985 35207 29019
rect 35207 28985 35216 29019
rect 35164 28976 35216 28985
rect 35808 28976 35860 29028
rect 35900 28976 35952 29028
rect 35992 28976 36044 29028
rect 39120 28976 39172 29028
rect 40776 29044 40828 29096
rect 31668 28951 31720 28960
rect 31668 28917 31677 28951
rect 31677 28917 31711 28951
rect 31711 28917 31720 28951
rect 31668 28908 31720 28917
rect 35256 28908 35308 28960
rect 35716 28908 35768 28960
rect 36084 28908 36136 28960
rect 37832 28908 37884 28960
rect 40040 28908 40092 28960
rect 42984 29112 43036 29164
rect 44088 29180 44140 29232
rect 46204 29180 46256 29232
rect 49884 29248 49936 29300
rect 43904 29112 43956 29164
rect 43812 29044 43864 29096
rect 44272 29087 44324 29096
rect 44272 29053 44281 29087
rect 44281 29053 44315 29087
rect 44315 29053 44324 29087
rect 44272 29044 44324 29053
rect 45100 29155 45152 29164
rect 45100 29121 45134 29155
rect 45134 29121 45152 29155
rect 45100 29112 45152 29121
rect 46112 29112 46164 29164
rect 46296 29112 46348 29164
rect 47676 29180 47728 29232
rect 46940 29155 46992 29164
rect 46940 29121 46949 29155
rect 46949 29121 46983 29155
rect 46983 29121 46992 29155
rect 46940 29112 46992 29121
rect 47492 29112 47544 29164
rect 47952 29155 48004 29164
rect 47952 29121 47959 29155
rect 47959 29121 48004 29155
rect 46480 29044 46532 29096
rect 46848 29044 46900 29096
rect 47952 29112 48004 29121
rect 48320 29112 48372 29164
rect 50160 29180 50212 29232
rect 55220 29248 55272 29300
rect 58348 29248 58400 29300
rect 54668 29180 54720 29232
rect 49516 29155 49568 29164
rect 49516 29121 49525 29155
rect 49525 29121 49559 29155
rect 49559 29121 49568 29155
rect 49700 29155 49752 29164
rect 49516 29112 49568 29121
rect 49700 29121 49709 29155
rect 49709 29121 49743 29155
rect 49743 29121 49752 29155
rect 49700 29112 49752 29121
rect 49884 29112 49936 29164
rect 50620 29112 50672 29164
rect 51356 29112 51408 29164
rect 51724 29112 51776 29164
rect 52828 29112 52880 29164
rect 53472 29112 53524 29164
rect 54392 29112 54444 29164
rect 55588 29180 55640 29232
rect 56692 29180 56744 29232
rect 53104 29044 53156 29096
rect 55404 29155 55456 29164
rect 55404 29121 55413 29155
rect 55413 29121 55447 29155
rect 55447 29121 55456 29155
rect 55404 29112 55456 29121
rect 55496 29155 55548 29164
rect 55496 29121 55505 29155
rect 55505 29121 55539 29155
rect 55539 29121 55548 29155
rect 55956 29155 56008 29164
rect 55496 29112 55548 29121
rect 55956 29121 55965 29155
rect 55965 29121 55999 29155
rect 55999 29121 56008 29155
rect 55956 29112 56008 29121
rect 56140 29112 56192 29164
rect 57336 29155 57388 29164
rect 44732 29019 44784 29028
rect 41604 28908 41656 28960
rect 44732 28985 44741 29019
rect 44741 28985 44775 29019
rect 44775 28985 44784 29019
rect 44732 28976 44784 28985
rect 47860 28976 47912 29028
rect 48136 28976 48188 29028
rect 57336 29121 57345 29155
rect 57345 29121 57379 29155
rect 57379 29121 57388 29155
rect 57336 29112 57388 29121
rect 42708 28951 42760 28960
rect 42708 28917 42717 28951
rect 42717 28917 42751 28951
rect 42751 28917 42760 28951
rect 42708 28908 42760 28917
rect 47032 28908 47084 28960
rect 48780 28908 48832 28960
rect 49148 28908 49200 28960
rect 49332 28908 49384 28960
rect 50804 28908 50856 28960
rect 51540 28951 51592 28960
rect 51540 28917 51549 28951
rect 51549 28917 51583 28951
rect 51583 28917 51592 28951
rect 51540 28908 51592 28917
rect 53472 28908 53524 28960
rect 53656 28951 53708 28960
rect 53656 28917 53665 28951
rect 53665 28917 53699 28951
rect 53699 28917 53708 28951
rect 53656 28908 53708 28917
rect 54852 28908 54904 28960
rect 55588 28908 55640 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 31208 28704 31260 28756
rect 34336 28747 34388 28756
rect 34336 28713 34345 28747
rect 34345 28713 34379 28747
rect 34379 28713 34388 28747
rect 34336 28704 34388 28713
rect 34612 28704 34664 28756
rect 34796 28704 34848 28756
rect 36912 28704 36964 28756
rect 37280 28704 37332 28756
rect 40040 28747 40092 28756
rect 40040 28713 40049 28747
rect 40049 28713 40083 28747
rect 40083 28713 40092 28747
rect 40040 28704 40092 28713
rect 40224 28704 40276 28756
rect 45192 28747 45244 28756
rect 36360 28636 36412 28688
rect 32312 28568 32364 28620
rect 33692 28568 33744 28620
rect 35808 28568 35860 28620
rect 38568 28636 38620 28688
rect 39672 28636 39724 28688
rect 32864 28500 32916 28552
rect 34796 28500 34848 28552
rect 35440 28500 35492 28552
rect 35900 28543 35952 28552
rect 35900 28509 35909 28543
rect 35909 28509 35943 28543
rect 35943 28509 35952 28543
rect 35900 28500 35952 28509
rect 35992 28543 36044 28552
rect 35992 28509 36001 28543
rect 36001 28509 36035 28543
rect 36035 28509 36044 28543
rect 37188 28568 37240 28620
rect 38384 28568 38436 28620
rect 35992 28500 36044 28509
rect 37556 28500 37608 28552
rect 38108 28543 38160 28552
rect 38108 28509 38117 28543
rect 38117 28509 38151 28543
rect 38151 28509 38160 28543
rect 38108 28500 38160 28509
rect 38200 28543 38252 28552
rect 38200 28509 38209 28543
rect 38209 28509 38243 28543
rect 38243 28509 38252 28543
rect 38200 28500 38252 28509
rect 38568 28500 38620 28552
rect 39948 28500 40000 28552
rect 40132 28543 40184 28552
rect 40132 28509 40141 28543
rect 40141 28509 40175 28543
rect 40175 28509 40184 28543
rect 40132 28500 40184 28509
rect 41144 28500 41196 28552
rect 42708 28568 42760 28620
rect 31668 28432 31720 28484
rect 33784 28432 33836 28484
rect 33140 28407 33192 28416
rect 33140 28373 33149 28407
rect 33149 28373 33183 28407
rect 33183 28373 33192 28407
rect 33140 28364 33192 28373
rect 35716 28364 35768 28416
rect 36084 28475 36136 28484
rect 36084 28441 36093 28475
rect 36093 28441 36127 28475
rect 36127 28441 36136 28475
rect 36084 28432 36136 28441
rect 37924 28432 37976 28484
rect 37372 28364 37424 28416
rect 38660 28364 38712 28416
rect 38936 28475 38988 28484
rect 38936 28441 38945 28475
rect 38945 28441 38979 28475
rect 38979 28441 38988 28475
rect 38936 28432 38988 28441
rect 39212 28432 39264 28484
rect 40868 28432 40920 28484
rect 41420 28475 41472 28484
rect 41420 28441 41429 28475
rect 41429 28441 41463 28475
rect 41463 28441 41472 28475
rect 41788 28500 41840 28552
rect 41420 28432 41472 28441
rect 41880 28432 41932 28484
rect 43260 28543 43312 28552
rect 43260 28509 43269 28543
rect 43269 28509 43303 28543
rect 43303 28509 43312 28543
rect 43260 28500 43312 28509
rect 45192 28713 45201 28747
rect 45201 28713 45235 28747
rect 45235 28713 45244 28747
rect 45192 28704 45244 28713
rect 45284 28704 45336 28756
rect 47676 28704 47728 28756
rect 44732 28636 44784 28688
rect 47308 28636 47360 28688
rect 48136 28636 48188 28688
rect 49332 28704 49384 28756
rect 49700 28704 49752 28756
rect 48872 28636 48924 28688
rect 50436 28636 50488 28688
rect 45192 28568 45244 28620
rect 45652 28543 45704 28552
rect 45652 28509 45697 28543
rect 45697 28509 45704 28543
rect 45652 28500 45704 28509
rect 45836 28543 45888 28552
rect 45836 28509 45845 28543
rect 45845 28509 45879 28543
rect 45879 28509 45888 28543
rect 46296 28543 46348 28552
rect 45836 28500 45888 28509
rect 46296 28509 46305 28543
rect 46305 28509 46339 28543
rect 46339 28509 46348 28543
rect 46296 28500 46348 28509
rect 46848 28568 46900 28620
rect 46664 28500 46716 28552
rect 48596 28568 48648 28620
rect 49148 28611 49200 28620
rect 49148 28577 49157 28611
rect 49157 28577 49191 28611
rect 49191 28577 49200 28611
rect 49148 28568 49200 28577
rect 52460 28704 52512 28756
rect 50804 28636 50856 28688
rect 54392 28679 54444 28688
rect 54392 28645 54401 28679
rect 54401 28645 54435 28679
rect 54435 28645 54444 28679
rect 54392 28636 54444 28645
rect 57336 28636 57388 28688
rect 54852 28611 54904 28620
rect 47492 28543 47544 28552
rect 47492 28509 47501 28543
rect 47501 28509 47535 28543
rect 47535 28509 47544 28543
rect 47492 28500 47544 28509
rect 47676 28500 47728 28552
rect 48228 28543 48280 28552
rect 48228 28509 48237 28543
rect 48237 28509 48271 28543
rect 48271 28509 48280 28543
rect 48228 28500 48280 28509
rect 49056 28543 49108 28552
rect 45192 28432 45244 28484
rect 47308 28432 47360 28484
rect 49056 28509 49065 28543
rect 49065 28509 49099 28543
rect 49099 28509 49108 28543
rect 49056 28500 49108 28509
rect 49424 28543 49476 28552
rect 49424 28509 49433 28543
rect 49433 28509 49467 28543
rect 49467 28509 49476 28543
rect 49424 28500 49476 28509
rect 50344 28543 50396 28552
rect 50344 28509 50353 28543
rect 50353 28509 50387 28543
rect 50387 28509 50396 28543
rect 50344 28500 50396 28509
rect 50528 28543 50580 28552
rect 50528 28509 50537 28543
rect 50537 28509 50571 28543
rect 50571 28509 50580 28543
rect 50528 28500 50580 28509
rect 50620 28500 50672 28552
rect 54852 28577 54861 28611
rect 54861 28577 54895 28611
rect 54895 28577 54904 28611
rect 54852 28568 54904 28577
rect 57520 28568 57572 28620
rect 51540 28500 51592 28552
rect 52276 28543 52328 28552
rect 52276 28509 52285 28543
rect 52285 28509 52319 28543
rect 52319 28509 52328 28543
rect 52276 28500 52328 28509
rect 53380 28543 53432 28552
rect 53380 28509 53389 28543
rect 53389 28509 53423 28543
rect 53423 28509 53432 28543
rect 53380 28500 53432 28509
rect 53472 28543 53524 28552
rect 53472 28509 53481 28543
rect 53481 28509 53515 28543
rect 53515 28509 53524 28543
rect 53472 28500 53524 28509
rect 53656 28543 53708 28552
rect 53656 28509 53691 28543
rect 53691 28509 53708 28543
rect 53656 28500 53708 28509
rect 54116 28500 54168 28552
rect 54760 28543 54812 28552
rect 54760 28509 54769 28543
rect 54769 28509 54803 28543
rect 54803 28509 54812 28543
rect 54760 28500 54812 28509
rect 57244 28500 57296 28552
rect 54024 28432 54076 28484
rect 41052 28407 41104 28416
rect 41052 28373 41061 28407
rect 41061 28373 41095 28407
rect 41095 28373 41104 28407
rect 41052 28364 41104 28373
rect 42156 28407 42208 28416
rect 42156 28373 42165 28407
rect 42165 28373 42199 28407
rect 42199 28373 42208 28407
rect 42156 28364 42208 28373
rect 42248 28364 42300 28416
rect 44272 28364 44324 28416
rect 46112 28364 46164 28416
rect 46756 28407 46808 28416
rect 46756 28373 46765 28407
rect 46765 28373 46799 28407
rect 46799 28373 46808 28407
rect 46756 28364 46808 28373
rect 47860 28364 47912 28416
rect 49332 28364 49384 28416
rect 51080 28407 51132 28416
rect 51080 28373 51089 28407
rect 51089 28373 51123 28407
rect 51123 28373 51132 28407
rect 51080 28364 51132 28373
rect 53932 28364 53984 28416
rect 56600 28407 56652 28416
rect 56600 28373 56609 28407
rect 56609 28373 56643 28407
rect 56643 28373 56652 28407
rect 56600 28364 56652 28373
rect 57244 28364 57296 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 37372 28160 37424 28212
rect 38292 28203 38344 28212
rect 38292 28169 38301 28203
rect 38301 28169 38335 28203
rect 38335 28169 38344 28203
rect 38292 28160 38344 28169
rect 40316 28160 40368 28212
rect 41788 28203 41840 28212
rect 33140 28092 33192 28144
rect 34336 28135 34388 28144
rect 34336 28101 34345 28135
rect 34345 28101 34379 28135
rect 34379 28101 34388 28135
rect 34336 28092 34388 28101
rect 34520 28092 34572 28144
rect 37556 28024 37608 28076
rect 39212 28024 39264 28076
rect 41788 28169 41797 28203
rect 41797 28169 41831 28203
rect 41831 28169 41840 28203
rect 41788 28160 41840 28169
rect 41880 28160 41932 28212
rect 43168 28160 43220 28212
rect 43720 28160 43772 28212
rect 44180 28160 44232 28212
rect 45468 28160 45520 28212
rect 46296 28160 46348 28212
rect 47124 28160 47176 28212
rect 49608 28160 49660 28212
rect 49700 28160 49752 28212
rect 50528 28160 50580 28212
rect 52000 28203 52052 28212
rect 32312 27999 32364 28008
rect 32312 27965 32321 27999
rect 32321 27965 32355 27999
rect 32355 27965 32364 27999
rect 32312 27956 32364 27965
rect 32588 27999 32640 28008
rect 32588 27965 32597 27999
rect 32597 27965 32631 27999
rect 32631 27965 32640 27999
rect 32588 27956 32640 27965
rect 38384 27956 38436 28008
rect 38568 27999 38620 28008
rect 38568 27965 38577 27999
rect 38577 27965 38611 27999
rect 38611 27965 38620 27999
rect 38568 27956 38620 27965
rect 39488 27956 39540 28008
rect 37280 27888 37332 27940
rect 42248 28024 42300 28076
rect 42524 28024 42576 28076
rect 31760 27863 31812 27872
rect 31760 27829 31769 27863
rect 31769 27829 31803 27863
rect 31803 27829 31812 27863
rect 31760 27820 31812 27829
rect 32956 27820 33008 27872
rect 39028 27820 39080 27872
rect 39488 27820 39540 27872
rect 40132 27956 40184 28008
rect 41972 27956 42024 28008
rect 43812 27956 43864 28008
rect 43996 28067 44048 28076
rect 43996 28033 44006 28067
rect 44006 28033 44040 28067
rect 44040 28033 44048 28067
rect 45284 28092 45336 28144
rect 43996 28024 44048 28033
rect 44272 28067 44324 28076
rect 44272 28033 44281 28067
rect 44281 28033 44315 28067
rect 44315 28033 44324 28067
rect 44272 28024 44324 28033
rect 45652 28024 45704 28076
rect 46388 28067 46440 28076
rect 45008 27956 45060 28008
rect 41420 27888 41472 27940
rect 45284 27999 45336 28008
rect 45284 27965 45293 27999
rect 45293 27965 45327 27999
rect 45327 27965 45336 27999
rect 45284 27956 45336 27965
rect 45928 27956 45980 28008
rect 46388 28033 46397 28067
rect 46397 28033 46431 28067
rect 46431 28033 46440 28067
rect 46388 28024 46440 28033
rect 46480 28067 46532 28076
rect 46480 28033 46489 28067
rect 46489 28033 46523 28067
rect 46523 28033 46532 28067
rect 46480 28024 46532 28033
rect 46664 28024 46716 28076
rect 47860 28024 47912 28076
rect 48044 28024 48096 28076
rect 48780 28067 48832 28076
rect 48780 28033 48789 28067
rect 48789 28033 48823 28067
rect 48823 28033 48832 28067
rect 48780 28024 48832 28033
rect 48964 28067 49016 28076
rect 48964 28033 48973 28067
rect 48973 28033 49007 28067
rect 49007 28033 49016 28067
rect 48964 28024 49016 28033
rect 50344 28092 50396 28144
rect 52000 28169 52009 28203
rect 52009 28169 52043 28203
rect 52043 28169 52052 28203
rect 52000 28160 52052 28169
rect 53380 28160 53432 28212
rect 55220 28160 55272 28212
rect 50620 28024 50672 28076
rect 52276 28092 52328 28144
rect 52828 28092 52880 28144
rect 53564 28092 53616 28144
rect 54024 28092 54076 28144
rect 51356 28067 51408 28076
rect 51356 28033 51365 28067
rect 51365 28033 51399 28067
rect 51399 28033 51408 28067
rect 51356 28024 51408 28033
rect 51540 28067 51592 28076
rect 51540 28033 51549 28067
rect 51549 28033 51583 28067
rect 51583 28033 51592 28067
rect 51540 28024 51592 28033
rect 54392 28067 54444 28076
rect 54392 28033 54401 28067
rect 54401 28033 54435 28067
rect 54435 28033 54444 28067
rect 54392 28024 54444 28033
rect 57152 28067 57204 28076
rect 57152 28033 57161 28067
rect 57161 28033 57195 28067
rect 57195 28033 57204 28067
rect 57152 28024 57204 28033
rect 58348 28067 58400 28076
rect 58348 28033 58357 28067
rect 58357 28033 58391 28067
rect 58391 28033 58400 28067
rect 58348 28024 58400 28033
rect 49608 27956 49660 28008
rect 40132 27820 40184 27872
rect 42984 27820 43036 27872
rect 45376 27820 45428 27872
rect 50252 27999 50304 28008
rect 50252 27965 50261 27999
rect 50261 27965 50295 27999
rect 50295 27965 50304 27999
rect 50252 27956 50304 27965
rect 50436 27956 50488 28008
rect 55588 27999 55640 28008
rect 54116 27931 54168 27940
rect 54116 27897 54125 27931
rect 54125 27897 54159 27931
rect 54159 27897 54168 27931
rect 54116 27888 54168 27897
rect 55588 27965 55597 27999
rect 55597 27965 55631 27999
rect 55631 27965 55640 27999
rect 55588 27956 55640 27965
rect 57244 27999 57296 28008
rect 57244 27965 57253 27999
rect 57253 27965 57287 27999
rect 57287 27965 57296 27999
rect 57244 27956 57296 27965
rect 58072 27999 58124 28008
rect 58072 27965 58081 27999
rect 58081 27965 58115 27999
rect 58115 27965 58124 27999
rect 58072 27956 58124 27965
rect 57336 27888 57388 27940
rect 47124 27820 47176 27872
rect 47952 27820 48004 27872
rect 49792 27820 49844 27872
rect 50528 27820 50580 27872
rect 51172 27820 51224 27872
rect 55864 27863 55916 27872
rect 55864 27829 55873 27863
rect 55873 27829 55907 27863
rect 55907 27829 55916 27863
rect 55864 27820 55916 27829
rect 56324 27863 56376 27872
rect 56324 27829 56333 27863
rect 56333 27829 56367 27863
rect 56367 27829 56376 27863
rect 56324 27820 56376 27829
rect 57704 27820 57756 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 32588 27659 32640 27668
rect 32588 27625 32597 27659
rect 32597 27625 32631 27659
rect 32631 27625 32640 27659
rect 32588 27616 32640 27625
rect 37188 27616 37240 27668
rect 38200 27616 38252 27668
rect 38568 27659 38620 27668
rect 38568 27625 38577 27659
rect 38577 27625 38611 27659
rect 38611 27625 38620 27659
rect 38568 27616 38620 27625
rect 39948 27616 40000 27668
rect 40132 27616 40184 27668
rect 40868 27616 40920 27668
rect 42156 27616 42208 27668
rect 43260 27616 43312 27668
rect 44364 27616 44416 27668
rect 45284 27616 45336 27668
rect 46388 27616 46440 27668
rect 47124 27616 47176 27668
rect 47676 27616 47728 27668
rect 36636 27548 36688 27600
rect 37280 27591 37332 27600
rect 37280 27557 37289 27591
rect 37289 27557 37323 27591
rect 37323 27557 37332 27591
rect 37280 27548 37332 27557
rect 33784 27455 33836 27464
rect 33784 27421 33793 27455
rect 33793 27421 33827 27455
rect 33827 27421 33836 27455
rect 33784 27412 33836 27421
rect 34612 27412 34664 27464
rect 36268 27480 36320 27532
rect 38752 27591 38804 27600
rect 38752 27557 38761 27591
rect 38761 27557 38795 27591
rect 38795 27557 38804 27591
rect 38752 27548 38804 27557
rect 39580 27548 39632 27600
rect 40592 27548 40644 27600
rect 46848 27548 46900 27600
rect 39028 27480 39080 27532
rect 38200 27455 38252 27464
rect 38200 27421 38209 27455
rect 38209 27421 38243 27455
rect 38243 27421 38252 27455
rect 38200 27412 38252 27421
rect 38660 27412 38712 27464
rect 39488 27455 39540 27464
rect 39488 27421 39497 27455
rect 39497 27421 39531 27455
rect 39531 27421 39540 27455
rect 39488 27412 39540 27421
rect 40684 27412 40736 27464
rect 41604 27480 41656 27532
rect 42708 27480 42760 27532
rect 44088 27455 44140 27464
rect 44088 27421 44097 27455
rect 44097 27421 44131 27455
rect 44131 27421 44140 27455
rect 44088 27412 44140 27421
rect 45376 27455 45428 27464
rect 45376 27421 45385 27455
rect 45385 27421 45419 27455
rect 45419 27421 45428 27455
rect 45376 27412 45428 27421
rect 45468 27412 45520 27464
rect 46112 27455 46164 27464
rect 46112 27421 46121 27455
rect 46121 27421 46155 27455
rect 46155 27421 46164 27455
rect 46112 27412 46164 27421
rect 46756 27412 46808 27464
rect 48044 27480 48096 27532
rect 47860 27455 47912 27464
rect 47860 27421 47869 27455
rect 47869 27421 47903 27455
rect 47903 27421 47912 27455
rect 47860 27412 47912 27421
rect 48136 27412 48188 27464
rect 49884 27616 49936 27668
rect 50436 27616 50488 27668
rect 51356 27616 51408 27668
rect 51540 27616 51592 27668
rect 53104 27616 53156 27668
rect 58072 27616 58124 27668
rect 48872 27548 48924 27600
rect 49608 27548 49660 27600
rect 53012 27591 53064 27600
rect 49516 27480 49568 27532
rect 51908 27523 51960 27532
rect 51908 27489 51917 27523
rect 51917 27489 51951 27523
rect 51951 27489 51960 27523
rect 51908 27480 51960 27489
rect 49608 27412 49660 27464
rect 50436 27412 50488 27464
rect 50620 27412 50672 27464
rect 51632 27455 51684 27464
rect 51632 27421 51641 27455
rect 51641 27421 51675 27455
rect 51675 27421 51684 27455
rect 51632 27412 51684 27421
rect 53012 27557 53021 27591
rect 53021 27557 53055 27591
rect 53055 27557 53064 27591
rect 53012 27548 53064 27557
rect 53104 27523 53156 27532
rect 53104 27489 53113 27523
rect 53113 27489 53147 27523
rect 53147 27489 53156 27523
rect 53104 27480 53156 27489
rect 53472 27480 53524 27532
rect 57796 27548 57848 27600
rect 36636 27344 36688 27396
rect 39212 27387 39264 27396
rect 33416 27276 33468 27328
rect 38476 27276 38528 27328
rect 39212 27353 39221 27387
rect 39221 27353 39255 27387
rect 39255 27353 39264 27387
rect 39212 27344 39264 27353
rect 42248 27344 42300 27396
rect 42984 27344 43036 27396
rect 41512 27276 41564 27328
rect 43904 27319 43956 27328
rect 43904 27285 43913 27319
rect 43913 27285 43947 27319
rect 43947 27285 43956 27319
rect 43904 27276 43956 27285
rect 44824 27276 44876 27328
rect 47952 27344 48004 27396
rect 47308 27276 47360 27328
rect 47492 27276 47544 27328
rect 48596 27344 48648 27396
rect 51264 27344 51316 27396
rect 49792 27276 49844 27328
rect 50896 27276 50948 27328
rect 52368 27276 52420 27328
rect 52736 27455 52788 27464
rect 52736 27421 52745 27455
rect 52745 27421 52779 27455
rect 52779 27421 52788 27455
rect 53932 27455 53984 27464
rect 52736 27412 52788 27421
rect 53932 27421 53941 27455
rect 53941 27421 53975 27455
rect 53975 27421 53984 27455
rect 53932 27412 53984 27421
rect 54300 27412 54352 27464
rect 54852 27412 54904 27464
rect 57704 27523 57756 27532
rect 57704 27489 57713 27523
rect 57713 27489 57747 27523
rect 57747 27489 57756 27523
rect 57704 27480 57756 27489
rect 55864 27455 55916 27464
rect 55864 27421 55873 27455
rect 55873 27421 55907 27455
rect 55907 27421 55916 27455
rect 55864 27412 55916 27421
rect 56508 27412 56560 27464
rect 56876 27344 56928 27396
rect 58072 27412 58124 27464
rect 58348 27412 58400 27464
rect 58164 27344 58216 27396
rect 54760 27276 54812 27328
rect 55036 27276 55088 27328
rect 55128 27276 55180 27328
rect 58256 27319 58308 27328
rect 58256 27285 58265 27319
rect 58265 27285 58299 27319
rect 58299 27285 58308 27319
rect 58256 27276 58308 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 33784 27072 33836 27124
rect 33416 27047 33468 27056
rect 33416 27013 33425 27047
rect 33425 27013 33459 27047
rect 33459 27013 33468 27047
rect 33416 27004 33468 27013
rect 34152 27004 34204 27056
rect 35348 27004 35400 27056
rect 39028 27115 39080 27124
rect 39028 27081 39037 27115
rect 39037 27081 39071 27115
rect 39071 27081 39080 27115
rect 39028 27072 39080 27081
rect 41328 27072 41380 27124
rect 45560 27115 45612 27124
rect 45560 27081 45569 27115
rect 45569 27081 45603 27115
rect 45603 27081 45612 27115
rect 45560 27072 45612 27081
rect 48044 27072 48096 27124
rect 37188 27004 37240 27056
rect 35992 26979 36044 26988
rect 35992 26945 36001 26979
rect 36001 26945 36035 26979
rect 36035 26945 36044 26979
rect 35992 26936 36044 26945
rect 40776 27004 40828 27056
rect 42524 27004 42576 27056
rect 43996 27004 44048 27056
rect 38476 26979 38528 26988
rect 32864 26732 32916 26784
rect 36268 26911 36320 26920
rect 36268 26877 36277 26911
rect 36277 26877 36311 26911
rect 36311 26877 36320 26911
rect 36268 26868 36320 26877
rect 37556 26843 37608 26852
rect 37556 26809 37565 26843
rect 37565 26809 37599 26843
rect 37599 26809 37608 26843
rect 37556 26800 37608 26809
rect 38476 26945 38485 26979
rect 38485 26945 38519 26979
rect 38519 26945 38528 26979
rect 38476 26936 38528 26945
rect 39488 26979 39540 26988
rect 39488 26945 39497 26979
rect 39497 26945 39531 26979
rect 39531 26945 39540 26979
rect 39488 26936 39540 26945
rect 39948 26936 40000 26988
rect 40684 26979 40736 26988
rect 40684 26945 40693 26979
rect 40693 26945 40727 26979
rect 40727 26945 40736 26979
rect 40684 26936 40736 26945
rect 41144 26979 41196 26988
rect 41144 26945 41153 26979
rect 41153 26945 41187 26979
rect 41187 26945 41196 26979
rect 41144 26936 41196 26945
rect 42984 26936 43036 26988
rect 37740 26868 37792 26920
rect 38200 26868 38252 26920
rect 40224 26868 40276 26920
rect 42432 26868 42484 26920
rect 44456 26936 44508 26988
rect 45100 27004 45152 27056
rect 45652 27004 45704 27056
rect 44824 26979 44876 26988
rect 44824 26945 44833 26979
rect 44833 26945 44867 26979
rect 44867 26945 44876 26979
rect 44824 26936 44876 26945
rect 45744 26936 45796 26988
rect 46296 26936 46348 26988
rect 46664 27004 46716 27056
rect 51264 27004 51316 27056
rect 46848 26936 46900 26988
rect 45836 26868 45888 26920
rect 46756 26868 46808 26920
rect 47676 26936 47728 26988
rect 48136 26936 48188 26988
rect 48964 26979 49016 26988
rect 48964 26945 48973 26979
rect 48973 26945 49007 26979
rect 49007 26945 49016 26979
rect 50068 26979 50120 26988
rect 48964 26936 49016 26945
rect 50068 26945 50077 26979
rect 50077 26945 50111 26979
rect 50111 26945 50120 26979
rect 50068 26936 50120 26945
rect 50160 26979 50212 26988
rect 50160 26945 50169 26979
rect 50169 26945 50203 26979
rect 50203 26945 50212 26979
rect 50344 26979 50396 26988
rect 50160 26936 50212 26945
rect 50344 26945 50353 26979
rect 50353 26945 50387 26979
rect 50387 26945 50396 26979
rect 50344 26936 50396 26945
rect 48872 26868 48924 26920
rect 49056 26868 49108 26920
rect 50528 26979 50580 26988
rect 50528 26945 50537 26979
rect 50537 26945 50571 26979
rect 50571 26945 50580 26979
rect 50528 26936 50580 26945
rect 51172 26936 51224 26988
rect 50896 26868 50948 26920
rect 54484 27072 54536 27124
rect 54760 27115 54812 27124
rect 54760 27081 54769 27115
rect 54769 27081 54803 27115
rect 54803 27081 54812 27115
rect 54760 27072 54812 27081
rect 52368 26936 52420 26988
rect 53196 27004 53248 27056
rect 55036 27047 55088 27056
rect 55036 27013 55045 27047
rect 55045 27013 55079 27047
rect 55079 27013 55088 27047
rect 55036 27004 55088 27013
rect 55128 27047 55180 27056
rect 55128 27013 55137 27047
rect 55137 27013 55171 27047
rect 55171 27013 55180 27047
rect 56876 27072 56928 27124
rect 55128 27004 55180 27013
rect 55864 27004 55916 27056
rect 53564 26936 53616 26988
rect 54668 26936 54720 26988
rect 56692 27004 56744 27056
rect 57888 27004 57940 27056
rect 53288 26911 53340 26920
rect 34612 26732 34664 26784
rect 38568 26775 38620 26784
rect 38568 26741 38577 26775
rect 38577 26741 38611 26775
rect 38611 26741 38620 26775
rect 38568 26732 38620 26741
rect 46388 26800 46440 26852
rect 46572 26800 46624 26852
rect 53288 26877 53297 26911
rect 53297 26877 53331 26911
rect 53331 26877 53340 26911
rect 53288 26868 53340 26877
rect 54300 26800 54352 26852
rect 43628 26732 43680 26784
rect 47032 26732 47084 26784
rect 48136 26732 48188 26784
rect 49608 26732 49660 26784
rect 51264 26732 51316 26784
rect 51632 26775 51684 26784
rect 51632 26741 51641 26775
rect 51641 26741 51675 26775
rect 51675 26741 51684 26775
rect 51632 26732 51684 26741
rect 52184 26775 52236 26784
rect 52184 26741 52193 26775
rect 52193 26741 52227 26775
rect 52227 26741 52236 26775
rect 52184 26732 52236 26741
rect 53472 26732 53524 26784
rect 53564 26732 53616 26784
rect 56600 26732 56652 26784
rect 58072 26775 58124 26784
rect 58072 26741 58081 26775
rect 58081 26741 58115 26775
rect 58115 26741 58124 26775
rect 58072 26732 58124 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2412 26528 2464 26580
rect 32312 26528 32364 26580
rect 32864 26528 32916 26580
rect 34152 26528 34204 26580
rect 36636 26571 36688 26580
rect 36636 26537 36645 26571
rect 36645 26537 36679 26571
rect 36679 26537 36688 26571
rect 36636 26528 36688 26537
rect 38936 26528 38988 26580
rect 39488 26528 39540 26580
rect 34704 26392 34756 26444
rect 40132 26460 40184 26512
rect 44088 26528 44140 26580
rect 45836 26528 45888 26580
rect 46848 26528 46900 26580
rect 42432 26503 42484 26512
rect 42432 26469 42441 26503
rect 42441 26469 42475 26503
rect 42475 26469 42484 26503
rect 42432 26460 42484 26469
rect 36452 26392 36504 26444
rect 38568 26392 38620 26444
rect 39212 26435 39264 26444
rect 39212 26401 39221 26435
rect 39221 26401 39255 26435
rect 39255 26401 39264 26435
rect 39212 26392 39264 26401
rect 40224 26392 40276 26444
rect 40316 26435 40368 26444
rect 40316 26401 40325 26435
rect 40325 26401 40359 26435
rect 40359 26401 40368 26435
rect 40316 26392 40368 26401
rect 41144 26392 41196 26444
rect 41328 26435 41380 26444
rect 41328 26401 41337 26435
rect 41337 26401 41371 26435
rect 41371 26401 41380 26435
rect 41328 26392 41380 26401
rect 32956 26367 33008 26376
rect 32956 26333 32965 26367
rect 32965 26333 32999 26367
rect 32999 26333 33008 26367
rect 32956 26324 33008 26333
rect 34796 26324 34848 26376
rect 37648 26367 37700 26376
rect 37648 26333 37657 26367
rect 37657 26333 37691 26367
rect 37691 26333 37700 26367
rect 37648 26324 37700 26333
rect 35164 26299 35216 26308
rect 35164 26265 35173 26299
rect 35173 26265 35207 26299
rect 35207 26265 35216 26299
rect 35164 26256 35216 26265
rect 36176 26256 36228 26308
rect 36544 26256 36596 26308
rect 37188 26256 37240 26308
rect 39672 26324 39724 26376
rect 40500 26324 40552 26376
rect 40684 26324 40736 26376
rect 41512 26324 41564 26376
rect 42708 26392 42760 26444
rect 45008 26324 45060 26376
rect 47216 26460 47268 26512
rect 47676 26460 47728 26512
rect 48872 26460 48924 26512
rect 46480 26435 46532 26444
rect 46480 26401 46489 26435
rect 46489 26401 46523 26435
rect 46523 26401 46532 26435
rect 46480 26392 46532 26401
rect 46756 26392 46808 26444
rect 47124 26324 47176 26376
rect 35992 26188 36044 26240
rect 38016 26188 38068 26240
rect 40316 26188 40368 26240
rect 43628 26256 43680 26308
rect 43904 26299 43956 26308
rect 43904 26265 43913 26299
rect 43913 26265 43947 26299
rect 43947 26265 43956 26299
rect 43904 26256 43956 26265
rect 45928 26256 45980 26308
rect 47492 26324 47544 26376
rect 48228 26392 48280 26444
rect 50620 26528 50672 26580
rect 52368 26571 52420 26580
rect 52368 26537 52377 26571
rect 52377 26537 52411 26571
rect 52411 26537 52420 26571
rect 52368 26528 52420 26537
rect 52920 26571 52972 26580
rect 52920 26537 52929 26571
rect 52929 26537 52963 26571
rect 52963 26537 52972 26571
rect 52920 26528 52972 26537
rect 53564 26571 53616 26580
rect 53564 26537 53573 26571
rect 53573 26537 53607 26571
rect 53607 26537 53616 26571
rect 53564 26528 53616 26537
rect 54300 26571 54352 26580
rect 54300 26537 54309 26571
rect 54309 26537 54343 26571
rect 54343 26537 54352 26571
rect 54300 26528 54352 26537
rect 54668 26571 54720 26580
rect 54668 26537 54677 26571
rect 54677 26537 54711 26571
rect 54711 26537 54720 26571
rect 54668 26528 54720 26537
rect 56324 26528 56376 26580
rect 56692 26571 56744 26580
rect 56692 26537 56701 26571
rect 56701 26537 56735 26571
rect 56735 26537 56744 26571
rect 56692 26528 56744 26537
rect 54484 26460 54536 26512
rect 48136 26324 48188 26376
rect 47676 26256 47728 26308
rect 48320 26256 48372 26308
rect 48964 26324 49016 26376
rect 49332 26367 49384 26376
rect 49332 26333 49341 26367
rect 49341 26333 49375 26367
rect 49375 26333 49384 26367
rect 49332 26324 49384 26333
rect 49700 26392 49752 26444
rect 54852 26392 54904 26444
rect 48780 26256 48832 26308
rect 49608 26324 49660 26376
rect 50528 26367 50580 26376
rect 50528 26333 50537 26367
rect 50537 26333 50571 26367
rect 50571 26333 50580 26367
rect 50528 26324 50580 26333
rect 51080 26324 51132 26376
rect 51264 26367 51316 26376
rect 51264 26333 51298 26367
rect 51298 26333 51316 26367
rect 51264 26324 51316 26333
rect 52276 26324 52328 26376
rect 51172 26256 51224 26308
rect 45836 26231 45888 26240
rect 45836 26197 45845 26231
rect 45845 26197 45879 26231
rect 45879 26197 45888 26231
rect 45836 26188 45888 26197
rect 46388 26188 46440 26240
rect 50528 26188 50580 26240
rect 50988 26188 51040 26240
rect 58072 26256 58124 26308
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 34704 25984 34756 26036
rect 35164 26027 35216 26036
rect 35164 25993 35173 26027
rect 35173 25993 35207 26027
rect 35207 25993 35216 26027
rect 35164 25984 35216 25993
rect 36268 25984 36320 26036
rect 39120 25984 39172 26036
rect 41420 25984 41472 26036
rect 42248 25984 42300 26036
rect 42616 25984 42668 26036
rect 43628 26027 43680 26036
rect 36636 25916 36688 25968
rect 37464 25848 37516 25900
rect 38016 25916 38068 25968
rect 41236 25916 41288 25968
rect 43628 25993 43637 26027
rect 43637 25993 43671 26027
rect 43671 25993 43680 26027
rect 43628 25984 43680 25993
rect 46296 26027 46348 26036
rect 46296 25993 46305 26027
rect 46305 25993 46339 26027
rect 46339 25993 46348 26027
rect 46296 25984 46348 25993
rect 46940 26027 46992 26036
rect 46940 25993 46949 26027
rect 46949 25993 46983 26027
rect 46983 25993 46992 26027
rect 46940 25984 46992 25993
rect 34796 25644 34848 25696
rect 35992 25780 36044 25832
rect 38016 25780 38068 25832
rect 38108 25644 38160 25696
rect 38660 25848 38712 25900
rect 40224 25848 40276 25900
rect 40500 25848 40552 25900
rect 41144 25848 41196 25900
rect 41972 25891 42024 25900
rect 41972 25857 41981 25891
rect 41981 25857 42015 25891
rect 42015 25857 42024 25891
rect 41972 25848 42024 25857
rect 42984 25848 43036 25900
rect 43996 25848 44048 25900
rect 45836 25848 45888 25900
rect 46020 25848 46072 25900
rect 47124 25916 47176 25968
rect 47584 25916 47636 25968
rect 49516 25984 49568 26036
rect 50988 25984 51040 26036
rect 52368 25984 52420 26036
rect 54576 26027 54628 26036
rect 54576 25993 54585 26027
rect 54585 25993 54619 26027
rect 54619 25993 54628 26027
rect 54576 25984 54628 25993
rect 56140 25984 56192 26036
rect 58256 25984 58308 26036
rect 47032 25848 47084 25900
rect 48228 25848 48280 25900
rect 39856 25780 39908 25832
rect 45928 25823 45980 25832
rect 45928 25789 45937 25823
rect 45937 25789 45971 25823
rect 45971 25789 45980 25823
rect 45928 25780 45980 25789
rect 48412 25891 48464 25900
rect 48412 25857 48421 25891
rect 48421 25857 48455 25891
rect 48455 25857 48464 25891
rect 50160 25916 50212 25968
rect 50804 25916 50856 25968
rect 48412 25848 48464 25857
rect 49792 25848 49844 25900
rect 49884 25891 49936 25900
rect 49884 25857 49893 25891
rect 49893 25857 49927 25891
rect 49927 25857 49936 25891
rect 49884 25848 49936 25857
rect 40040 25712 40092 25764
rect 47860 25712 47912 25764
rect 50804 25712 50856 25764
rect 38936 25644 38988 25696
rect 44180 25644 44232 25696
rect 44364 25644 44416 25696
rect 44916 25687 44968 25696
rect 44916 25653 44925 25687
rect 44925 25653 44959 25687
rect 44959 25653 44968 25687
rect 44916 25644 44968 25653
rect 48688 25644 48740 25696
rect 48872 25687 48924 25696
rect 48872 25653 48881 25687
rect 48881 25653 48915 25687
rect 48915 25653 48924 25687
rect 48872 25644 48924 25653
rect 51540 25687 51592 25696
rect 51540 25653 51549 25687
rect 51549 25653 51583 25687
rect 51583 25653 51592 25687
rect 51540 25644 51592 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 36176 25440 36228 25492
rect 37464 25483 37516 25492
rect 37464 25449 37473 25483
rect 37473 25449 37507 25483
rect 37507 25449 37516 25483
rect 37464 25440 37516 25449
rect 38016 25483 38068 25492
rect 38016 25449 38025 25483
rect 38025 25449 38059 25483
rect 38059 25449 38068 25483
rect 38016 25440 38068 25449
rect 38108 25440 38160 25492
rect 39120 25483 39172 25492
rect 39120 25449 39129 25483
rect 39129 25449 39163 25483
rect 39163 25449 39172 25483
rect 39120 25440 39172 25449
rect 40132 25440 40184 25492
rect 40500 25483 40552 25492
rect 40500 25449 40509 25483
rect 40509 25449 40543 25483
rect 40543 25449 40552 25483
rect 40500 25440 40552 25449
rect 41144 25440 41196 25492
rect 43076 25440 43128 25492
rect 43812 25440 43864 25492
rect 46296 25440 46348 25492
rect 47308 25440 47360 25492
rect 48228 25483 48280 25492
rect 48228 25449 48237 25483
rect 48237 25449 48271 25483
rect 48271 25449 48280 25483
rect 48228 25440 48280 25449
rect 49056 25483 49108 25492
rect 49056 25449 49065 25483
rect 49065 25449 49099 25483
rect 49099 25449 49108 25483
rect 49056 25440 49108 25449
rect 37648 25304 37700 25356
rect 39856 25372 39908 25424
rect 31760 25236 31812 25288
rect 36452 25279 36504 25288
rect 34796 25100 34848 25152
rect 36452 25245 36461 25279
rect 36461 25245 36495 25279
rect 36495 25245 36504 25279
rect 36452 25236 36504 25245
rect 37004 25236 37056 25288
rect 38200 25279 38252 25288
rect 36544 25168 36596 25220
rect 38200 25245 38209 25279
rect 38209 25245 38243 25279
rect 38243 25245 38252 25279
rect 38200 25236 38252 25245
rect 38476 25279 38528 25288
rect 38476 25245 38485 25279
rect 38485 25245 38519 25279
rect 38519 25245 38528 25279
rect 38476 25236 38528 25245
rect 39028 25279 39080 25288
rect 39028 25245 39037 25279
rect 39037 25245 39071 25279
rect 39071 25245 39080 25279
rect 39028 25236 39080 25245
rect 38844 25168 38896 25220
rect 40408 25304 40460 25356
rect 40868 25304 40920 25356
rect 43168 25372 43220 25424
rect 46480 25372 46532 25424
rect 48412 25372 48464 25424
rect 52184 25440 52236 25492
rect 52644 25415 52696 25424
rect 42708 25304 42760 25356
rect 45100 25236 45152 25288
rect 46204 25236 46256 25288
rect 52644 25381 52653 25415
rect 52653 25381 52687 25415
rect 52687 25381 52696 25415
rect 52644 25372 52696 25381
rect 57980 25372 58032 25424
rect 49884 25304 49936 25356
rect 50068 25304 50120 25356
rect 47032 25279 47084 25288
rect 47032 25245 47041 25279
rect 47041 25245 47075 25279
rect 47075 25245 47084 25279
rect 47032 25236 47084 25245
rect 47216 25279 47268 25288
rect 47216 25245 47225 25279
rect 47225 25245 47259 25279
rect 47259 25245 47268 25279
rect 47216 25236 47268 25245
rect 47308 25279 47360 25288
rect 47308 25245 47317 25279
rect 47317 25245 47351 25279
rect 47351 25245 47360 25279
rect 48320 25279 48372 25288
rect 47308 25236 47360 25245
rect 48320 25245 48329 25279
rect 48329 25245 48363 25279
rect 48363 25245 48372 25279
rect 48320 25236 48372 25245
rect 39856 25100 39908 25152
rect 40316 25143 40368 25152
rect 40316 25109 40325 25143
rect 40325 25109 40359 25143
rect 40359 25109 40368 25143
rect 40316 25100 40368 25109
rect 41052 25168 41104 25220
rect 43076 25168 43128 25220
rect 46940 25168 46992 25220
rect 49608 25236 49660 25288
rect 50160 25236 50212 25288
rect 51080 25304 51132 25356
rect 50988 25236 51040 25288
rect 51816 25236 51868 25288
rect 42248 25100 42300 25152
rect 45192 25100 45244 25152
rect 46296 25143 46348 25152
rect 46296 25109 46305 25143
rect 46305 25109 46339 25143
rect 46339 25109 46348 25143
rect 46296 25100 46348 25109
rect 47584 25100 47636 25152
rect 48228 25100 48280 25152
rect 49700 25168 49752 25220
rect 51080 25168 51132 25220
rect 51632 25100 51684 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 36452 24896 36504 24948
rect 37556 24896 37608 24948
rect 34612 24803 34664 24812
rect 34612 24769 34621 24803
rect 34621 24769 34655 24803
rect 34655 24769 34664 24803
rect 34612 24760 34664 24769
rect 35992 24760 36044 24812
rect 37464 24828 37516 24880
rect 38844 24871 38896 24880
rect 38844 24837 38853 24871
rect 38853 24837 38887 24871
rect 38887 24837 38896 24871
rect 38844 24828 38896 24837
rect 37832 24803 37884 24812
rect 37832 24769 37841 24803
rect 37841 24769 37875 24803
rect 37875 24769 37884 24803
rect 37832 24760 37884 24769
rect 38936 24803 38988 24812
rect 38936 24769 38945 24803
rect 38945 24769 38979 24803
rect 38979 24769 38988 24803
rect 38936 24760 38988 24769
rect 40132 24896 40184 24948
rect 40868 24896 40920 24948
rect 40040 24871 40092 24880
rect 39396 24760 39448 24812
rect 40040 24837 40049 24871
rect 40049 24837 40083 24871
rect 40083 24837 40092 24871
rect 40040 24828 40092 24837
rect 40316 24828 40368 24880
rect 41604 24828 41656 24880
rect 38844 24692 38896 24744
rect 38292 24624 38344 24676
rect 39672 24667 39724 24676
rect 39672 24633 39681 24667
rect 39681 24633 39715 24667
rect 39715 24633 39724 24667
rect 39672 24624 39724 24633
rect 40408 24760 40460 24812
rect 40868 24803 40920 24812
rect 40868 24769 40877 24803
rect 40877 24769 40911 24803
rect 40911 24769 40920 24803
rect 40868 24760 40920 24769
rect 40960 24760 41012 24812
rect 39948 24692 40000 24744
rect 41788 24735 41840 24744
rect 41788 24701 41797 24735
rect 41797 24701 41831 24735
rect 41831 24701 41840 24735
rect 41788 24692 41840 24701
rect 45928 24828 45980 24880
rect 41972 24760 42024 24812
rect 42892 24803 42944 24812
rect 42892 24769 42901 24803
rect 42901 24769 42935 24803
rect 42935 24769 42944 24803
rect 42892 24760 42944 24769
rect 45192 24760 45244 24812
rect 45376 24760 45428 24812
rect 46940 24760 46992 24812
rect 47860 24803 47912 24812
rect 47860 24769 47869 24803
rect 47869 24769 47903 24803
rect 47903 24769 47912 24803
rect 47860 24760 47912 24769
rect 48780 24803 48832 24812
rect 48780 24769 48789 24803
rect 48789 24769 48823 24803
rect 48823 24769 48832 24803
rect 48780 24760 48832 24769
rect 51172 24803 51224 24812
rect 51172 24769 51181 24803
rect 51181 24769 51215 24803
rect 51215 24769 51224 24803
rect 51172 24760 51224 24769
rect 42708 24692 42760 24744
rect 44180 24692 44232 24744
rect 51080 24692 51132 24744
rect 37556 24556 37608 24608
rect 39028 24556 39080 24608
rect 39304 24556 39356 24608
rect 39856 24599 39908 24608
rect 39856 24565 39865 24599
rect 39865 24565 39899 24599
rect 39899 24565 39908 24599
rect 39856 24556 39908 24565
rect 41052 24667 41104 24676
rect 41052 24633 41061 24667
rect 41061 24633 41095 24667
rect 41095 24633 41104 24667
rect 41052 24624 41104 24633
rect 41604 24599 41656 24608
rect 41604 24565 41613 24599
rect 41613 24565 41647 24599
rect 41647 24565 41656 24599
rect 47032 24624 47084 24676
rect 48688 24624 48740 24676
rect 52644 24760 52696 24812
rect 51632 24692 51684 24744
rect 41604 24556 41656 24565
rect 47584 24556 47636 24608
rect 50252 24599 50304 24608
rect 50252 24565 50261 24599
rect 50261 24565 50295 24599
rect 50295 24565 50304 24599
rect 50252 24556 50304 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 35992 24352 36044 24404
rect 40776 24352 40828 24404
rect 43076 24352 43128 24404
rect 44916 24352 44968 24404
rect 47032 24352 47084 24404
rect 48320 24352 48372 24404
rect 50344 24352 50396 24404
rect 37372 24284 37424 24336
rect 38476 24284 38528 24336
rect 37188 24259 37240 24268
rect 37188 24225 37197 24259
rect 37197 24225 37231 24259
rect 37231 24225 37240 24259
rect 37188 24216 37240 24225
rect 38016 24259 38068 24268
rect 38016 24225 38025 24259
rect 38025 24225 38059 24259
rect 38059 24225 38068 24259
rect 40040 24284 40092 24336
rect 45376 24284 45428 24336
rect 38016 24216 38068 24225
rect 35992 24148 36044 24200
rect 38292 24191 38344 24200
rect 38292 24157 38301 24191
rect 38301 24157 38335 24191
rect 38335 24157 38344 24191
rect 39028 24191 39080 24200
rect 38292 24148 38344 24157
rect 39028 24157 39037 24191
rect 39037 24157 39071 24191
rect 39071 24157 39080 24191
rect 39028 24148 39080 24157
rect 40960 24216 41012 24268
rect 46296 24259 46348 24268
rect 46296 24225 46305 24259
rect 46305 24225 46339 24259
rect 46339 24225 46348 24259
rect 46296 24216 46348 24225
rect 47676 24259 47728 24268
rect 47676 24225 47685 24259
rect 47685 24225 47719 24259
rect 47719 24225 47728 24259
rect 47676 24216 47728 24225
rect 49608 24216 49660 24268
rect 39764 24148 39816 24200
rect 39856 24148 39908 24200
rect 40868 24191 40920 24200
rect 40868 24157 40877 24191
rect 40877 24157 40911 24191
rect 40911 24157 40920 24191
rect 40868 24148 40920 24157
rect 37832 24080 37884 24132
rect 35072 24055 35124 24064
rect 35072 24021 35081 24055
rect 35081 24021 35115 24055
rect 35115 24021 35124 24055
rect 35072 24012 35124 24021
rect 38844 24055 38896 24064
rect 38844 24021 38853 24055
rect 38853 24021 38887 24055
rect 38887 24021 38896 24055
rect 38844 24012 38896 24021
rect 40316 24080 40368 24132
rect 41604 24191 41656 24200
rect 41604 24157 41613 24191
rect 41613 24157 41647 24191
rect 41647 24157 41656 24191
rect 41604 24148 41656 24157
rect 40500 24012 40552 24064
rect 42156 24080 42208 24132
rect 42892 24148 42944 24200
rect 43444 24148 43496 24200
rect 45100 24148 45152 24200
rect 47400 24191 47452 24200
rect 46204 24080 46256 24132
rect 47400 24157 47409 24191
rect 47409 24157 47443 24191
rect 47443 24157 47452 24191
rect 47400 24148 47452 24157
rect 49700 24148 49752 24200
rect 51080 24148 51132 24200
rect 45284 24055 45336 24064
rect 45284 24021 45293 24055
rect 45293 24021 45327 24055
rect 45327 24021 45336 24055
rect 45284 24012 45336 24021
rect 46296 24055 46348 24064
rect 46296 24021 46305 24055
rect 46305 24021 46339 24055
rect 46339 24021 46348 24055
rect 46296 24012 46348 24021
rect 49056 24080 49108 24132
rect 49884 24012 49936 24064
rect 51448 24055 51500 24064
rect 51448 24021 51457 24055
rect 51457 24021 51491 24055
rect 51491 24021 51500 24055
rect 51448 24012 51500 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 34704 23808 34756 23860
rect 36544 23851 36596 23860
rect 36544 23817 36553 23851
rect 36553 23817 36587 23851
rect 36587 23817 36596 23851
rect 36544 23808 36596 23817
rect 37188 23808 37240 23860
rect 37832 23808 37884 23860
rect 39764 23851 39816 23860
rect 39764 23817 39773 23851
rect 39773 23817 39807 23851
rect 39807 23817 39816 23851
rect 39764 23808 39816 23817
rect 40316 23851 40368 23860
rect 40316 23817 40325 23851
rect 40325 23817 40359 23851
rect 40359 23817 40368 23851
rect 40316 23808 40368 23817
rect 35072 23783 35124 23792
rect 35072 23749 35081 23783
rect 35081 23749 35115 23783
rect 35115 23749 35124 23783
rect 35072 23740 35124 23749
rect 36084 23740 36136 23792
rect 38384 23740 38436 23792
rect 40776 23808 40828 23860
rect 41052 23808 41104 23860
rect 41328 23740 41380 23792
rect 46296 23808 46348 23860
rect 46388 23808 46440 23860
rect 49056 23808 49108 23860
rect 38016 23672 38068 23724
rect 39856 23672 39908 23724
rect 42064 23715 42116 23724
rect 42064 23681 42073 23715
rect 42073 23681 42107 23715
rect 42107 23681 42116 23715
rect 42064 23672 42116 23681
rect 42708 23672 42760 23724
rect 45284 23740 45336 23792
rect 46020 23783 46072 23792
rect 46020 23749 46029 23783
rect 46029 23749 46063 23783
rect 46063 23749 46072 23783
rect 46020 23740 46072 23749
rect 49792 23783 49844 23792
rect 49792 23749 49801 23783
rect 49801 23749 49835 23783
rect 49835 23749 49844 23783
rect 49792 23740 49844 23749
rect 51448 23740 51500 23792
rect 43444 23715 43496 23724
rect 43444 23681 43453 23715
rect 43453 23681 43487 23715
rect 43487 23681 43496 23715
rect 43444 23672 43496 23681
rect 46940 23672 46992 23724
rect 47768 23715 47820 23724
rect 47768 23681 47777 23715
rect 47777 23681 47811 23715
rect 47811 23681 47820 23715
rect 47768 23672 47820 23681
rect 48780 23672 48832 23724
rect 49148 23672 49200 23724
rect 51816 23715 51868 23724
rect 51816 23681 51825 23715
rect 51825 23681 51859 23715
rect 51859 23681 51868 23715
rect 51816 23672 51868 23681
rect 35440 23604 35492 23656
rect 49884 23604 49936 23656
rect 38476 23468 38528 23520
rect 41328 23468 41380 23520
rect 42984 23468 43036 23520
rect 47032 23536 47084 23588
rect 46848 23468 46900 23520
rect 49148 23468 49200 23520
rect 51080 23468 51132 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 35440 23264 35492 23316
rect 38108 23264 38160 23316
rect 41788 23264 41840 23316
rect 46940 23264 46992 23316
rect 51816 23307 51868 23316
rect 51816 23273 51825 23307
rect 51825 23273 51859 23307
rect 51859 23273 51868 23307
rect 51816 23264 51868 23273
rect 36084 23196 36136 23248
rect 37832 23128 37884 23180
rect 35992 23060 36044 23112
rect 37188 23103 37240 23112
rect 37188 23069 37197 23103
rect 37197 23069 37231 23103
rect 37231 23069 37240 23103
rect 37188 23060 37240 23069
rect 37372 23103 37424 23112
rect 37372 23069 37381 23103
rect 37381 23069 37415 23103
rect 37415 23069 37424 23103
rect 37372 23060 37424 23069
rect 39856 23128 39908 23180
rect 42064 23128 42116 23180
rect 38844 23060 38896 23112
rect 39396 23103 39448 23112
rect 39396 23069 39405 23103
rect 39405 23069 39439 23103
rect 39439 23069 39448 23103
rect 39396 23060 39448 23069
rect 42984 23103 43036 23112
rect 42984 23069 42993 23103
rect 42993 23069 43027 23103
rect 43027 23069 43036 23103
rect 42984 23060 43036 23069
rect 49884 23196 49936 23248
rect 47216 23128 47268 23180
rect 48872 23171 48924 23180
rect 48872 23137 48881 23171
rect 48881 23137 48915 23171
rect 48915 23137 48924 23171
rect 48872 23128 48924 23137
rect 37648 22992 37700 23044
rect 39212 22992 39264 23044
rect 40776 22992 40828 23044
rect 42156 22992 42208 23044
rect 42800 22992 42852 23044
rect 43444 22992 43496 23044
rect 49792 23060 49844 23112
rect 50252 23060 50304 23112
rect 46204 22992 46256 23044
rect 46480 23035 46532 23044
rect 46480 23001 46489 23035
rect 46489 23001 46523 23035
rect 46523 23001 46532 23035
rect 46480 22992 46532 23001
rect 47124 22992 47176 23044
rect 37280 22924 37332 22976
rect 38200 22924 38252 22976
rect 38568 22924 38620 22976
rect 39304 22967 39356 22976
rect 39304 22933 39313 22967
rect 39313 22933 39347 22967
rect 39347 22933 39356 22967
rect 39304 22924 39356 22933
rect 43904 22967 43956 22976
rect 43904 22933 43913 22967
rect 43913 22933 43947 22967
rect 43947 22933 43956 22967
rect 43904 22924 43956 22933
rect 44456 22924 44508 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 37556 22763 37608 22772
rect 37556 22729 37565 22763
rect 37565 22729 37599 22763
rect 37599 22729 37608 22763
rect 37556 22720 37608 22729
rect 39856 22763 39908 22772
rect 39856 22729 39865 22763
rect 39865 22729 39899 22763
rect 39899 22729 39908 22763
rect 39856 22720 39908 22729
rect 40776 22763 40828 22772
rect 40776 22729 40785 22763
rect 40785 22729 40819 22763
rect 40819 22729 40828 22763
rect 40776 22720 40828 22729
rect 41512 22720 41564 22772
rect 43904 22720 43956 22772
rect 37372 22584 37424 22636
rect 38016 22652 38068 22704
rect 39120 22652 39172 22704
rect 38108 22627 38160 22636
rect 38108 22593 38117 22627
rect 38117 22593 38151 22627
rect 38151 22593 38160 22627
rect 38108 22584 38160 22593
rect 42800 22652 42852 22704
rect 44456 22695 44508 22704
rect 44456 22661 44465 22695
rect 44465 22661 44499 22695
rect 44499 22661 44508 22695
rect 44456 22652 44508 22661
rect 46480 22720 46532 22772
rect 49700 22720 49752 22772
rect 51080 22763 51132 22772
rect 51080 22729 51089 22763
rect 51089 22729 51123 22763
rect 51123 22729 51132 22763
rect 51080 22720 51132 22729
rect 46204 22695 46256 22704
rect 46204 22661 46213 22695
rect 46213 22661 46247 22695
rect 46247 22661 46256 22695
rect 46204 22652 46256 22661
rect 38384 22559 38436 22568
rect 38384 22525 38393 22559
rect 38393 22525 38427 22559
rect 38427 22525 38436 22559
rect 38384 22516 38436 22525
rect 36268 22423 36320 22432
rect 36268 22389 36277 22423
rect 36277 22389 36311 22423
rect 36311 22389 36320 22423
rect 36268 22380 36320 22389
rect 37648 22380 37700 22432
rect 42708 22584 42760 22636
rect 46848 22627 46900 22636
rect 46848 22593 46857 22627
rect 46857 22593 46891 22627
rect 46891 22593 46900 22627
rect 46848 22584 46900 22593
rect 47400 22584 47452 22636
rect 49424 22584 49476 22636
rect 48320 22559 48372 22568
rect 48320 22525 48329 22559
rect 48329 22525 48363 22559
rect 48363 22525 48372 22559
rect 48320 22516 48372 22525
rect 51540 22380 51592 22432
rect 58164 22380 58216 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 36268 22219 36320 22228
rect 36268 22185 36298 22219
rect 36298 22185 36320 22219
rect 36268 22176 36320 22185
rect 48320 22176 48372 22228
rect 37372 22108 37424 22160
rect 35440 22083 35492 22092
rect 35440 22049 35449 22083
rect 35449 22049 35483 22083
rect 35483 22049 35492 22083
rect 35440 22040 35492 22049
rect 39212 22040 39264 22092
rect 47124 22040 47176 22092
rect 38476 22015 38528 22024
rect 38476 21981 38485 22015
rect 38485 21981 38519 22015
rect 38519 21981 38528 22015
rect 38476 21972 38528 21981
rect 38752 21972 38804 22024
rect 37556 21904 37608 21956
rect 38568 21904 38620 21956
rect 47032 21972 47084 22024
rect 48228 22040 48280 22092
rect 49148 22040 49200 22092
rect 49424 22040 49476 22092
rect 38660 21836 38712 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 37556 21675 37608 21684
rect 37556 21641 37565 21675
rect 37565 21641 37599 21675
rect 37599 21641 37608 21675
rect 37556 21632 37608 21641
rect 38384 21632 38436 21684
rect 39120 21632 39172 21684
rect 47768 21675 47820 21684
rect 47768 21641 47777 21675
rect 47777 21641 47811 21675
rect 47811 21641 47820 21675
rect 47768 21632 47820 21641
rect 37648 21539 37700 21548
rect 37648 21505 37657 21539
rect 37657 21505 37691 21539
rect 37691 21505 37700 21539
rect 37648 21496 37700 21505
rect 38660 21496 38712 21548
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 47308 21131 47360 21140
rect 47308 21097 47317 21131
rect 47317 21097 47351 21131
rect 47351 21097 47360 21131
rect 47308 21088 47360 21097
rect 50344 20884 50396 20936
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 58624 2796 58676 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 1952 2592 2004 2644
rect 34704 2592 34756 2644
rect 58164 2635 58216 2644
rect 58164 2601 58173 2635
rect 58173 2601 58207 2635
rect 58207 2601 58216 2635
rect 58164 2592 58216 2601
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 29000 2252 29052 2304
rect 58624 2320 58676 2372
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
rect 20 1300 72 1352
rect 1584 1300 1636 1352
<< metal2 >>
rect 1306 59200 1362 59800
rect 30930 59200 30986 59800
rect 59910 59200 59966 59800
rect 1320 57458 1348 59200
rect 4874 57692 5182 57701
rect 4874 57690 4880 57692
rect 4936 57690 4960 57692
rect 5016 57690 5040 57692
rect 5096 57690 5120 57692
rect 5176 57690 5182 57692
rect 4936 57638 4938 57690
rect 5118 57638 5120 57690
rect 4874 57636 4880 57638
rect 4936 57636 4960 57638
rect 5016 57636 5040 57638
rect 5096 57636 5120 57638
rect 5176 57636 5182 57638
rect 4874 57627 5182 57636
rect 1308 57452 1360 57458
rect 1308 57394 1360 57400
rect 1952 57248 2004 57254
rect 1952 57190 2004 57196
rect 2044 57248 2096 57254
rect 2044 57190 2096 57196
rect 1964 56846 1992 57190
rect 1952 56840 2004 56846
rect 1952 56782 2004 56788
rect 2056 56710 2084 57190
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 2136 56908 2188 56914
rect 2136 56850 2188 56856
rect 1584 56704 1636 56710
rect 1584 56646 1636 56652
rect 2044 56704 2096 56710
rect 2044 56646 2096 56652
rect 1596 56438 1624 56646
rect 1584 56432 1636 56438
rect 1584 56374 1636 56380
rect 2056 56166 2084 56646
rect 2044 56160 2096 56166
rect 2044 56102 2096 56108
rect 2148 45554 2176 56850
rect 4874 56604 5182 56613
rect 4874 56602 4880 56604
rect 4936 56602 4960 56604
rect 5016 56602 5040 56604
rect 5096 56602 5120 56604
rect 5176 56602 5182 56604
rect 4936 56550 4938 56602
rect 5118 56550 5120 56602
rect 4874 56548 4880 56550
rect 4936 56548 4960 56550
rect 5016 56548 5040 56550
rect 5096 56548 5120 56550
rect 5176 56548 5182 56550
rect 4874 56539 5182 56548
rect 30944 56506 30972 59200
rect 35594 57692 35902 57701
rect 35594 57690 35600 57692
rect 35656 57690 35680 57692
rect 35736 57690 35760 57692
rect 35816 57690 35840 57692
rect 35896 57690 35902 57692
rect 35656 57638 35658 57690
rect 35838 57638 35840 57690
rect 35594 57636 35600 57638
rect 35656 57636 35680 57638
rect 35736 57636 35760 57638
rect 35816 57636 35840 57638
rect 35896 57636 35902 57638
rect 35594 57627 35902 57636
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 59924 56846 59952 59200
rect 58348 56840 58400 56846
rect 58348 56782 58400 56788
rect 59912 56840 59964 56846
rect 59912 56782 59964 56788
rect 35594 56604 35902 56613
rect 35594 56602 35600 56604
rect 35656 56602 35680 56604
rect 35736 56602 35760 56604
rect 35816 56602 35840 56604
rect 35896 56602 35902 56604
rect 35656 56550 35658 56602
rect 35838 56550 35840 56602
rect 35594 56548 35600 56550
rect 35656 56548 35680 56550
rect 35736 56548 35760 56550
rect 35816 56548 35840 56550
rect 35896 56548 35902 56550
rect 35594 56539 35902 56548
rect 58360 56506 58388 56782
rect 58624 56704 58676 56710
rect 58624 56646 58676 56652
rect 30380 56500 30432 56506
rect 30380 56442 30432 56448
rect 30932 56500 30984 56506
rect 30932 56442 30984 56448
rect 58348 56500 58400 56506
rect 58348 56442 58400 56448
rect 30392 56166 30420 56442
rect 30380 56160 30432 56166
rect 30380 56102 30432 56108
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4874 55516 5182 55525
rect 4874 55514 4880 55516
rect 4936 55514 4960 55516
rect 5016 55514 5040 55516
rect 5096 55514 5120 55516
rect 5176 55514 5182 55516
rect 4936 55462 4938 55514
rect 5118 55462 5120 55514
rect 4874 55460 4880 55462
rect 4936 55460 4960 55462
rect 5016 55460 5040 55462
rect 5096 55460 5120 55462
rect 5176 55460 5182 55462
rect 4874 55451 5182 55460
rect 30392 55214 30420 56102
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 35594 55516 35902 55525
rect 35594 55514 35600 55516
rect 35656 55514 35680 55516
rect 35736 55514 35760 55516
rect 35816 55514 35840 55516
rect 35896 55514 35902 55516
rect 35656 55462 35658 55514
rect 35838 55462 35840 55514
rect 35594 55460 35600 55462
rect 35656 55460 35680 55462
rect 35736 55460 35760 55462
rect 35816 55460 35840 55462
rect 35896 55460 35902 55462
rect 35594 55451 35902 55460
rect 30392 55186 30512 55214
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4874 54428 5182 54437
rect 4874 54426 4880 54428
rect 4936 54426 4960 54428
rect 5016 54426 5040 54428
rect 5096 54426 5120 54428
rect 5176 54426 5182 54428
rect 4936 54374 4938 54426
rect 5118 54374 5120 54426
rect 4874 54372 4880 54374
rect 4936 54372 4960 54374
rect 5016 54372 5040 54374
rect 5096 54372 5120 54374
rect 5176 54372 5182 54374
rect 4874 54363 5182 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4874 53340 5182 53349
rect 4874 53338 4880 53340
rect 4936 53338 4960 53340
rect 5016 53338 5040 53340
rect 5096 53338 5120 53340
rect 5176 53338 5182 53340
rect 4936 53286 4938 53338
rect 5118 53286 5120 53338
rect 4874 53284 4880 53286
rect 4936 53284 4960 53286
rect 5016 53284 5040 53286
rect 5096 53284 5120 53286
rect 5176 53284 5182 53286
rect 4874 53275 5182 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4874 52252 5182 52261
rect 4874 52250 4880 52252
rect 4936 52250 4960 52252
rect 5016 52250 5040 52252
rect 5096 52250 5120 52252
rect 5176 52250 5182 52252
rect 4936 52198 4938 52250
rect 5118 52198 5120 52250
rect 4874 52196 4880 52198
rect 4936 52196 4960 52198
rect 5016 52196 5040 52198
rect 5096 52196 5120 52198
rect 5176 52196 5182 52198
rect 4874 52187 5182 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4874 51164 5182 51173
rect 4874 51162 4880 51164
rect 4936 51162 4960 51164
rect 5016 51162 5040 51164
rect 5096 51162 5120 51164
rect 5176 51162 5182 51164
rect 4936 51110 4938 51162
rect 5118 51110 5120 51162
rect 4874 51108 4880 51110
rect 4936 51108 4960 51110
rect 5016 51108 5040 51110
rect 5096 51108 5120 51110
rect 5176 51108 5182 51110
rect 4874 51099 5182 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4874 50076 5182 50085
rect 4874 50074 4880 50076
rect 4936 50074 4960 50076
rect 5016 50074 5040 50076
rect 5096 50074 5120 50076
rect 5176 50074 5182 50076
rect 4936 50022 4938 50074
rect 5118 50022 5120 50074
rect 4874 50020 4880 50022
rect 4936 50020 4960 50022
rect 5016 50020 5040 50022
rect 5096 50020 5120 50022
rect 5176 50020 5182 50022
rect 4874 50011 5182 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4874 48988 5182 48997
rect 4874 48986 4880 48988
rect 4936 48986 4960 48988
rect 5016 48986 5040 48988
rect 5096 48986 5120 48988
rect 5176 48986 5182 48988
rect 4936 48934 4938 48986
rect 5118 48934 5120 48986
rect 4874 48932 4880 48934
rect 4936 48932 4960 48934
rect 5016 48932 5040 48934
rect 5096 48932 5120 48934
rect 5176 48932 5182 48934
rect 4874 48923 5182 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4874 47900 5182 47909
rect 4874 47898 4880 47900
rect 4936 47898 4960 47900
rect 5016 47898 5040 47900
rect 5096 47898 5120 47900
rect 5176 47898 5182 47900
rect 4936 47846 4938 47898
rect 5118 47846 5120 47898
rect 4874 47844 4880 47846
rect 4936 47844 4960 47846
rect 5016 47844 5040 47846
rect 5096 47844 5120 47846
rect 5176 47844 5182 47846
rect 4874 47835 5182 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4874 46812 5182 46821
rect 4874 46810 4880 46812
rect 4936 46810 4960 46812
rect 5016 46810 5040 46812
rect 5096 46810 5120 46812
rect 5176 46810 5182 46812
rect 4936 46758 4938 46810
rect 5118 46758 5120 46810
rect 4874 46756 4880 46758
rect 4936 46756 4960 46758
rect 5016 46756 5040 46758
rect 5096 46756 5120 46758
rect 5176 46756 5182 46758
rect 4874 46747 5182 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4874 45724 5182 45733
rect 4874 45722 4880 45724
rect 4936 45722 4960 45724
rect 5016 45722 5040 45724
rect 5096 45722 5120 45724
rect 5176 45722 5182 45724
rect 4936 45670 4938 45722
rect 5118 45670 5120 45722
rect 4874 45668 4880 45670
rect 4936 45668 4960 45670
rect 5016 45668 5040 45670
rect 5096 45668 5120 45670
rect 5176 45668 5182 45670
rect 4874 45659 5182 45668
rect 1964 45526 2176 45554
rect 1674 30696 1730 30705
rect 1674 30631 1730 30640
rect 1688 30598 1716 30631
rect 1676 30592 1728 30598
rect 1676 30534 1728 30540
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1596 2446 1624 2790
rect 1964 2650 1992 45526
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4874 44636 5182 44645
rect 4874 44634 4880 44636
rect 4936 44634 4960 44636
rect 5016 44634 5040 44636
rect 5096 44634 5120 44636
rect 5176 44634 5182 44636
rect 4936 44582 4938 44634
rect 5118 44582 5120 44634
rect 4874 44580 4880 44582
rect 4936 44580 4960 44582
rect 5016 44580 5040 44582
rect 5096 44580 5120 44582
rect 5176 44580 5182 44582
rect 4874 44571 5182 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 30012 43240 30064 43246
rect 30012 43182 30064 43188
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 30024 42226 30052 43182
rect 30196 42764 30248 42770
rect 30196 42706 30248 42712
rect 30012 42220 30064 42226
rect 30012 42162 30064 42168
rect 29276 42152 29328 42158
rect 29276 42094 29328 42100
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 28908 41676 28960 41682
rect 28908 41618 28960 41624
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 28920 40526 28948 41618
rect 29288 41614 29316 42094
rect 29276 41608 29328 41614
rect 29276 41550 29328 41556
rect 29092 41064 29144 41070
rect 29092 41006 29144 41012
rect 29104 40730 29132 41006
rect 29092 40724 29144 40730
rect 29092 40666 29144 40672
rect 28908 40520 28960 40526
rect 28908 40462 28960 40468
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 28816 37324 28868 37330
rect 28816 37266 28868 37272
rect 28172 37256 28224 37262
rect 28172 37198 28224 37204
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 28184 36786 28212 37198
rect 28264 37120 28316 37126
rect 28264 37062 28316 37068
rect 28276 36922 28304 37062
rect 28828 36938 28856 37266
rect 28920 37210 28948 40462
rect 29184 39976 29236 39982
rect 29184 39918 29236 39924
rect 29000 39840 29052 39846
rect 29000 39782 29052 39788
rect 29012 39642 29040 39782
rect 29000 39636 29052 39642
rect 29000 39578 29052 39584
rect 29196 39506 29224 39918
rect 29184 39500 29236 39506
rect 29184 39442 29236 39448
rect 29196 38894 29224 39442
rect 29184 38888 29236 38894
rect 29184 38830 29236 38836
rect 29288 38010 29316 41550
rect 29828 40588 29880 40594
rect 29828 40530 29880 40536
rect 29840 39438 29868 40530
rect 29828 39432 29880 39438
rect 29828 39374 29880 39380
rect 29736 38956 29788 38962
rect 29736 38898 29788 38904
rect 29748 38282 29776 38898
rect 29736 38276 29788 38282
rect 29736 38218 29788 38224
rect 29276 38004 29328 38010
rect 29276 37946 29328 37952
rect 29184 37868 29236 37874
rect 29184 37810 29236 37816
rect 28920 37182 29132 37210
rect 29104 37126 29132 37182
rect 28908 37120 28960 37126
rect 29092 37120 29144 37126
rect 28960 37068 29040 37074
rect 28908 37062 29040 37068
rect 29092 37062 29144 37068
rect 28920 37046 29040 37062
rect 29012 36938 29040 37046
rect 28264 36916 28316 36922
rect 28828 36910 28948 36938
rect 29012 36910 29132 36938
rect 28264 36858 28316 36864
rect 28172 36780 28224 36786
rect 28172 36722 28224 36728
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 27344 35012 27396 35018
rect 27344 34954 27396 34960
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 27356 34610 27384 34954
rect 27620 34740 27672 34746
rect 27620 34682 27672 34688
rect 27344 34604 27396 34610
rect 27344 34546 27396 34552
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 27632 33930 27660 34682
rect 28080 34536 28132 34542
rect 28080 34478 28132 34484
rect 28092 34202 28120 34478
rect 28080 34196 28132 34202
rect 28080 34138 28132 34144
rect 27620 33924 27672 33930
rect 27620 33866 27672 33872
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 28092 33522 28120 34138
rect 28080 33516 28132 33522
rect 28080 33458 28132 33464
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 28276 31482 28304 36858
rect 28920 36786 28948 36910
rect 29104 36786 29132 36910
rect 28908 36780 28960 36786
rect 28908 36722 28960 36728
rect 29092 36780 29144 36786
rect 29092 36722 29144 36728
rect 28920 36174 28948 36722
rect 29104 36530 29132 36722
rect 29196 36650 29224 37810
rect 29276 37664 29328 37670
rect 29276 37606 29328 37612
rect 29288 37194 29316 37606
rect 29368 37324 29420 37330
rect 29368 37266 29420 37272
rect 29276 37188 29328 37194
rect 29276 37130 29328 37136
rect 29288 36650 29316 37130
rect 29380 36718 29408 37266
rect 29748 36922 29776 38218
rect 29736 36916 29788 36922
rect 29736 36858 29788 36864
rect 29368 36712 29420 36718
rect 29368 36654 29420 36660
rect 29184 36644 29236 36650
rect 29184 36586 29236 36592
rect 29276 36644 29328 36650
rect 29276 36586 29328 36592
rect 29104 36502 29224 36530
rect 28908 36168 28960 36174
rect 28908 36110 28960 36116
rect 28356 36032 28408 36038
rect 28356 35974 28408 35980
rect 28368 32502 28396 35974
rect 28920 35766 28948 36110
rect 29196 36106 29224 36502
rect 29276 36168 29328 36174
rect 29276 36110 29328 36116
rect 29184 36100 29236 36106
rect 29184 36042 29236 36048
rect 28908 35760 28960 35766
rect 28908 35702 28960 35708
rect 28920 35154 28948 35702
rect 29196 35698 29224 36042
rect 29184 35692 29236 35698
rect 29184 35634 29236 35640
rect 29288 35562 29316 36110
rect 29276 35556 29328 35562
rect 29276 35498 29328 35504
rect 28908 35148 28960 35154
rect 28908 35090 28960 35096
rect 29000 35080 29052 35086
rect 29000 35022 29052 35028
rect 29012 34746 29040 35022
rect 29000 34740 29052 34746
rect 29000 34682 29052 34688
rect 29092 34672 29144 34678
rect 29092 34614 29144 34620
rect 28540 34400 28592 34406
rect 28540 34342 28592 34348
rect 28356 32496 28408 32502
rect 28356 32438 28408 32444
rect 28264 31476 28316 31482
rect 28264 31418 28316 31424
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 2412 30592 2464 30598
rect 2412 30534 2464 30540
rect 2424 26586 2452 30534
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 28552 30122 28580 34342
rect 29104 34202 29132 34614
rect 29092 34196 29144 34202
rect 29092 34138 29144 34144
rect 29184 33992 29236 33998
rect 29184 33934 29236 33940
rect 28908 33924 28960 33930
rect 28908 33866 28960 33872
rect 28920 30258 28948 33866
rect 29196 33318 29224 33934
rect 29184 33312 29236 33318
rect 29184 33254 29236 33260
rect 29196 33114 29224 33254
rect 29184 33108 29236 33114
rect 29184 33050 29236 33056
rect 29196 32910 29224 33050
rect 29184 32904 29236 32910
rect 29184 32846 29236 32852
rect 28816 30252 28868 30258
rect 28816 30194 28868 30200
rect 28908 30252 28960 30258
rect 28908 30194 28960 30200
rect 28540 30116 28592 30122
rect 28540 30058 28592 30064
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 28828 29510 28856 30194
rect 29380 29850 29408 36654
rect 29748 36122 29776 36858
rect 29840 36310 29868 39374
rect 30024 36922 30052 42162
rect 30208 42158 30236 42706
rect 30196 42152 30248 42158
rect 30196 42094 30248 42100
rect 30380 40452 30432 40458
rect 30380 40394 30432 40400
rect 30392 39982 30420 40394
rect 30380 39976 30432 39982
rect 30380 39918 30432 39924
rect 30392 39370 30420 39918
rect 30380 39364 30432 39370
rect 30380 39306 30432 39312
rect 30380 38752 30432 38758
rect 30380 38694 30432 38700
rect 30392 38350 30420 38694
rect 30104 38344 30156 38350
rect 30380 38344 30432 38350
rect 30156 38304 30236 38332
rect 30104 38286 30156 38292
rect 30208 37806 30236 38304
rect 30380 38286 30432 38292
rect 30380 37868 30432 37874
rect 30380 37810 30432 37816
rect 30196 37800 30248 37806
rect 30196 37742 30248 37748
rect 30208 37194 30236 37742
rect 30196 37188 30248 37194
rect 30196 37130 30248 37136
rect 30012 36916 30064 36922
rect 30012 36858 30064 36864
rect 30208 36854 30236 37130
rect 30196 36848 30248 36854
rect 30196 36790 30248 36796
rect 29920 36780 29972 36786
rect 29920 36722 29972 36728
rect 29932 36378 29960 36722
rect 29920 36372 29972 36378
rect 29920 36314 29972 36320
rect 29828 36304 29880 36310
rect 29828 36246 29880 36252
rect 29748 36106 29868 36122
rect 29748 36100 29880 36106
rect 29748 36094 29828 36100
rect 29828 36042 29880 36048
rect 29460 35828 29512 35834
rect 29460 35770 29512 35776
rect 29472 30802 29500 35770
rect 30104 35692 30156 35698
rect 30104 35634 30156 35640
rect 30116 35290 30144 35634
rect 30104 35284 30156 35290
rect 30104 35226 30156 35232
rect 30208 34678 30236 36790
rect 30392 36718 30420 37810
rect 30380 36712 30432 36718
rect 30380 36654 30432 36660
rect 30380 36236 30432 36242
rect 30380 36178 30432 36184
rect 30392 35850 30420 36178
rect 30300 35834 30420 35850
rect 30288 35828 30420 35834
rect 30340 35822 30420 35828
rect 30288 35770 30340 35776
rect 30484 34950 30512 55186
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 35594 54428 35902 54437
rect 35594 54426 35600 54428
rect 35656 54426 35680 54428
rect 35736 54426 35760 54428
rect 35816 54426 35840 54428
rect 35896 54426 35902 54428
rect 35656 54374 35658 54426
rect 35838 54374 35840 54426
rect 35594 54372 35600 54374
rect 35656 54372 35680 54374
rect 35736 54372 35760 54374
rect 35816 54372 35840 54374
rect 35896 54372 35902 54374
rect 35594 54363 35902 54372
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 35594 53340 35902 53349
rect 35594 53338 35600 53340
rect 35656 53338 35680 53340
rect 35736 53338 35760 53340
rect 35816 53338 35840 53340
rect 35896 53338 35902 53340
rect 35656 53286 35658 53338
rect 35838 53286 35840 53338
rect 35594 53284 35600 53286
rect 35656 53284 35680 53286
rect 35736 53284 35760 53286
rect 35816 53284 35840 53286
rect 35896 53284 35902 53286
rect 35594 53275 35902 53284
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 35594 52252 35902 52261
rect 35594 52250 35600 52252
rect 35656 52250 35680 52252
rect 35736 52250 35760 52252
rect 35816 52250 35840 52252
rect 35896 52250 35902 52252
rect 35656 52198 35658 52250
rect 35838 52198 35840 52250
rect 35594 52196 35600 52198
rect 35656 52196 35680 52198
rect 35736 52196 35760 52198
rect 35816 52196 35840 52198
rect 35896 52196 35902 52198
rect 35594 52187 35902 52196
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 35594 51164 35902 51173
rect 35594 51162 35600 51164
rect 35656 51162 35680 51164
rect 35736 51162 35760 51164
rect 35816 51162 35840 51164
rect 35896 51162 35902 51164
rect 35656 51110 35658 51162
rect 35838 51110 35840 51162
rect 35594 51108 35600 51110
rect 35656 51108 35680 51110
rect 35736 51108 35760 51110
rect 35816 51108 35840 51110
rect 35896 51108 35902 51110
rect 35594 51099 35902 51108
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 35594 50076 35902 50085
rect 35594 50074 35600 50076
rect 35656 50074 35680 50076
rect 35736 50074 35760 50076
rect 35816 50074 35840 50076
rect 35896 50074 35902 50076
rect 35656 50022 35658 50074
rect 35838 50022 35840 50074
rect 35594 50020 35600 50022
rect 35656 50020 35680 50022
rect 35736 50020 35760 50022
rect 35816 50020 35840 50022
rect 35896 50020 35902 50022
rect 35594 50011 35902 50020
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 35594 48988 35902 48997
rect 35594 48986 35600 48988
rect 35656 48986 35680 48988
rect 35736 48986 35760 48988
rect 35816 48986 35840 48988
rect 35896 48986 35902 48988
rect 35656 48934 35658 48986
rect 35838 48934 35840 48986
rect 35594 48932 35600 48934
rect 35656 48932 35680 48934
rect 35736 48932 35760 48934
rect 35816 48932 35840 48934
rect 35896 48932 35902 48934
rect 35594 48923 35902 48932
rect 43352 48816 43404 48822
rect 43352 48758 43404 48764
rect 35348 48748 35400 48754
rect 35348 48690 35400 48696
rect 37648 48748 37700 48754
rect 37648 48690 37700 48696
rect 40224 48748 40276 48754
rect 40224 48690 40276 48696
rect 40592 48748 40644 48754
rect 40592 48690 40644 48696
rect 40960 48748 41012 48754
rect 40960 48690 41012 48696
rect 42800 48748 42852 48754
rect 42852 48708 42932 48736
rect 42800 48690 42852 48696
rect 33140 48544 33192 48550
rect 33140 48486 33192 48492
rect 34244 48544 34296 48550
rect 34244 48486 34296 48492
rect 34796 48544 34848 48550
rect 34796 48486 34848 48492
rect 32588 48136 32640 48142
rect 32588 48078 32640 48084
rect 32496 47660 32548 47666
rect 32496 47602 32548 47608
rect 31668 47524 31720 47530
rect 31668 47466 31720 47472
rect 31484 45960 31536 45966
rect 31484 45902 31536 45908
rect 31496 45554 31524 45902
rect 31576 45554 31628 45558
rect 31496 45552 31628 45554
rect 31496 45526 31576 45552
rect 31116 45280 31168 45286
rect 31116 45222 31168 45228
rect 31128 44878 31156 45222
rect 31116 44872 31168 44878
rect 31116 44814 31168 44820
rect 31024 44328 31076 44334
rect 31024 44270 31076 44276
rect 31036 43314 31064 44270
rect 31116 43784 31168 43790
rect 31116 43726 31168 43732
rect 31024 43308 31076 43314
rect 31024 43250 31076 43256
rect 31036 41750 31064 43250
rect 31128 43246 31156 43726
rect 31116 43240 31168 43246
rect 31116 43182 31168 43188
rect 31392 42696 31444 42702
rect 31392 42638 31444 42644
rect 31116 42220 31168 42226
rect 31116 42162 31168 42168
rect 31024 41744 31076 41750
rect 31024 41686 31076 41692
rect 30656 41676 30708 41682
rect 30656 41618 30708 41624
rect 30668 41414 30696 41618
rect 30840 41608 30892 41614
rect 30840 41550 30892 41556
rect 30668 41386 30788 41414
rect 30564 40520 30616 40526
rect 30564 40462 30616 40468
rect 30576 39574 30604 40462
rect 30656 40044 30708 40050
rect 30656 39986 30708 39992
rect 30668 39642 30696 39986
rect 30656 39636 30708 39642
rect 30656 39578 30708 39584
rect 30564 39568 30616 39574
rect 30564 39510 30616 39516
rect 30656 39432 30708 39438
rect 30656 39374 30708 39380
rect 30564 39364 30616 39370
rect 30564 39306 30616 39312
rect 30576 39098 30604 39306
rect 30564 39092 30616 39098
rect 30564 39034 30616 39040
rect 30668 38554 30696 39374
rect 30656 38548 30708 38554
rect 30656 38490 30708 38496
rect 30760 38434 30788 41386
rect 30852 40730 30880 41550
rect 30840 40724 30892 40730
rect 30840 40666 30892 40672
rect 30840 40452 30892 40458
rect 30840 40394 30892 40400
rect 30932 40452 30984 40458
rect 30932 40394 30984 40400
rect 30852 40186 30880 40394
rect 30840 40180 30892 40186
rect 30840 40122 30892 40128
rect 30944 40050 30972 40394
rect 31128 40050 31156 42162
rect 30932 40044 30984 40050
rect 30932 39986 30984 39992
rect 31116 40044 31168 40050
rect 31116 39986 31168 39992
rect 30840 38956 30892 38962
rect 30840 38898 30892 38904
rect 30668 38406 30788 38434
rect 30564 37936 30616 37942
rect 30564 37878 30616 37884
rect 30576 37262 30604 37878
rect 30668 37466 30696 38406
rect 30748 38208 30800 38214
rect 30748 38150 30800 38156
rect 30656 37460 30708 37466
rect 30656 37402 30708 37408
rect 30760 37330 30788 38150
rect 30852 37806 30880 38898
rect 30932 37868 30984 37874
rect 30932 37810 30984 37816
rect 30840 37800 30892 37806
rect 30840 37742 30892 37748
rect 30944 37330 30972 37810
rect 30748 37324 30800 37330
rect 30748 37266 30800 37272
rect 30932 37324 30984 37330
rect 30932 37266 30984 37272
rect 30564 37256 30616 37262
rect 30564 37198 30616 37204
rect 30576 36786 30604 37198
rect 30944 36786 30972 37266
rect 30564 36780 30616 36786
rect 30564 36722 30616 36728
rect 30932 36780 30984 36786
rect 30932 36722 30984 36728
rect 30576 36174 30604 36722
rect 30656 36712 30708 36718
rect 30656 36654 30708 36660
rect 30564 36168 30616 36174
rect 30564 36110 30616 36116
rect 30576 35766 30604 36110
rect 30668 36038 30696 36654
rect 30944 36242 30972 36722
rect 30932 36236 30984 36242
rect 30932 36178 30984 36184
rect 30656 36032 30708 36038
rect 30656 35974 30708 35980
rect 30564 35760 30616 35766
rect 30564 35702 30616 35708
rect 30656 35080 30708 35086
rect 30656 35022 30708 35028
rect 30472 34944 30524 34950
rect 30472 34886 30524 34892
rect 30668 34678 30696 35022
rect 30196 34672 30248 34678
rect 30196 34614 30248 34620
rect 30656 34672 30708 34678
rect 30656 34614 30708 34620
rect 30668 34202 30696 34614
rect 30656 34196 30708 34202
rect 30656 34138 30708 34144
rect 29736 34060 29788 34066
rect 29736 34002 29788 34008
rect 29748 33522 29776 34002
rect 30564 33924 30616 33930
rect 30564 33866 30616 33872
rect 29736 33516 29788 33522
rect 29736 33458 29788 33464
rect 29748 32978 29776 33458
rect 30576 33114 30604 33866
rect 31024 33584 31076 33590
rect 31024 33526 31076 33532
rect 30564 33108 30616 33114
rect 30564 33050 30616 33056
rect 29736 32972 29788 32978
rect 29736 32914 29788 32920
rect 29644 32768 29696 32774
rect 29644 32710 29696 32716
rect 29656 32502 29684 32710
rect 29748 32570 29776 32914
rect 30288 32904 30340 32910
rect 30288 32846 30340 32852
rect 30300 32570 30328 32846
rect 31036 32570 31064 33526
rect 29736 32564 29788 32570
rect 29736 32506 29788 32512
rect 30288 32564 30340 32570
rect 30288 32506 30340 32512
rect 31024 32564 31076 32570
rect 31024 32506 31076 32512
rect 29644 32496 29696 32502
rect 29644 32438 29696 32444
rect 30196 32496 30248 32502
rect 30196 32438 30248 32444
rect 30208 31958 30236 32438
rect 30300 32026 30328 32506
rect 31128 32026 31156 39986
rect 31404 39914 31432 42638
rect 31392 39908 31444 39914
rect 31392 39850 31444 39856
rect 31392 39636 31444 39642
rect 31392 39578 31444 39584
rect 31404 39370 31432 39578
rect 31392 39364 31444 39370
rect 31392 39306 31444 39312
rect 31206 38584 31262 38593
rect 31206 38519 31262 38528
rect 31220 38350 31248 38519
rect 31208 38344 31260 38350
rect 31208 38286 31260 38292
rect 31208 37868 31260 37874
rect 31208 37810 31260 37816
rect 31220 35698 31248 37810
rect 31404 36854 31432 39306
rect 31496 38010 31524 45526
rect 31576 45494 31628 45500
rect 31680 44878 31708 47466
rect 32220 47184 32272 47190
rect 32220 47126 32272 47132
rect 32232 47054 32260 47126
rect 32220 47048 32272 47054
rect 32220 46990 32272 46996
rect 32128 46980 32180 46986
rect 32128 46922 32180 46928
rect 31760 46572 31812 46578
rect 31760 46514 31812 46520
rect 31772 46170 31800 46514
rect 31852 46368 31904 46374
rect 31852 46310 31904 46316
rect 31760 46164 31812 46170
rect 31760 46106 31812 46112
rect 31864 45830 31892 46310
rect 32140 45966 32168 46922
rect 32128 45960 32180 45966
rect 32128 45902 32180 45908
rect 31852 45824 31904 45830
rect 31852 45766 31904 45772
rect 31864 45626 31892 45766
rect 31852 45620 31904 45626
rect 31852 45562 31904 45568
rect 31852 45416 31904 45422
rect 31852 45358 31904 45364
rect 31864 44946 31892 45358
rect 31852 44940 31904 44946
rect 31852 44882 31904 44888
rect 31668 44872 31720 44878
rect 31668 44814 31720 44820
rect 31680 44402 31708 44814
rect 31668 44396 31720 44402
rect 31668 44338 31720 44344
rect 31864 42770 31892 44882
rect 32232 44198 32260 46990
rect 32312 46912 32364 46918
rect 32312 46854 32364 46860
rect 32324 45966 32352 46854
rect 32508 46170 32536 47602
rect 32600 47598 32628 48078
rect 33152 48006 33180 48486
rect 33140 48000 33192 48006
rect 33140 47942 33192 47948
rect 33152 47734 33180 47942
rect 33140 47728 33192 47734
rect 33140 47670 33192 47676
rect 32588 47592 32640 47598
rect 32588 47534 32640 47540
rect 32600 46714 32628 47534
rect 32864 47116 32916 47122
rect 32864 47058 32916 47064
rect 32680 47048 32732 47054
rect 32680 46990 32732 46996
rect 32588 46708 32640 46714
rect 32588 46650 32640 46656
rect 32692 46374 32720 46990
rect 32772 46436 32824 46442
rect 32772 46378 32824 46384
rect 32680 46368 32732 46374
rect 32680 46310 32732 46316
rect 32496 46164 32548 46170
rect 32496 46106 32548 46112
rect 32588 46096 32640 46102
rect 32508 46044 32588 46050
rect 32508 46038 32640 46044
rect 32508 46022 32628 46038
rect 32692 46034 32720 46310
rect 32680 46028 32732 46034
rect 32312 45960 32364 45966
rect 32312 45902 32364 45908
rect 32404 45824 32456 45830
rect 32404 45766 32456 45772
rect 32416 45490 32444 45766
rect 32404 45484 32456 45490
rect 32404 45426 32456 45432
rect 32416 44946 32444 45426
rect 32404 44940 32456 44946
rect 32404 44882 32456 44888
rect 32508 44742 32536 46022
rect 32680 45970 32732 45976
rect 32784 44878 32812 46378
rect 32876 44962 32904 47058
rect 33152 46918 33180 47670
rect 32956 46912 33008 46918
rect 32956 46854 33008 46860
rect 33140 46912 33192 46918
rect 33140 46854 33192 46860
rect 32968 45898 32996 46854
rect 34256 46646 34284 48486
rect 34704 48068 34756 48074
rect 34704 48010 34756 48016
rect 34520 47456 34572 47462
rect 34520 47398 34572 47404
rect 34532 46918 34560 47398
rect 34520 46912 34572 46918
rect 34520 46854 34572 46860
rect 34244 46640 34296 46646
rect 34244 46582 34296 46588
rect 33600 46572 33652 46578
rect 33600 46514 33652 46520
rect 33324 46504 33376 46510
rect 33324 46446 33376 46452
rect 33336 46034 33364 46446
rect 33612 46374 33640 46514
rect 33784 46504 33836 46510
rect 33784 46446 33836 46452
rect 33600 46368 33652 46374
rect 33600 46310 33652 46316
rect 33324 46028 33376 46034
rect 33324 45970 33376 45976
rect 32956 45892 33008 45898
rect 32956 45834 33008 45840
rect 32968 45801 32996 45834
rect 33048 45824 33100 45830
rect 32954 45792 33010 45801
rect 33048 45766 33100 45772
rect 32954 45727 33010 45736
rect 32876 44934 32996 44962
rect 32772 44872 32824 44878
rect 32772 44814 32824 44820
rect 32864 44872 32916 44878
rect 32864 44814 32916 44820
rect 32496 44736 32548 44742
rect 32496 44678 32548 44684
rect 32404 44328 32456 44334
rect 32404 44270 32456 44276
rect 32220 44192 32272 44198
rect 32220 44134 32272 44140
rect 31852 42764 31904 42770
rect 31852 42706 31904 42712
rect 31760 42696 31812 42702
rect 31760 42638 31812 42644
rect 32220 42696 32272 42702
rect 32220 42638 32272 42644
rect 31772 42362 31800 42638
rect 32232 42362 32260 42638
rect 31760 42356 31812 42362
rect 31760 42298 31812 42304
rect 32220 42356 32272 42362
rect 32220 42298 32272 42304
rect 32220 42220 32272 42226
rect 32220 42162 32272 42168
rect 31852 41676 31904 41682
rect 31852 41618 31904 41624
rect 31864 41041 31892 41618
rect 32232 41614 32260 42162
rect 32416 42090 32444 44270
rect 32508 42702 32536 44678
rect 32588 44192 32640 44198
rect 32588 44134 32640 44140
rect 32496 42696 32548 42702
rect 32600 42684 32628 44134
rect 32680 43784 32732 43790
rect 32680 43726 32732 43732
rect 32692 42838 32720 43726
rect 32680 42832 32732 42838
rect 32680 42774 32732 42780
rect 32600 42656 32720 42684
rect 32496 42638 32548 42644
rect 32404 42084 32456 42090
rect 32404 42026 32456 42032
rect 31944 41608 31996 41614
rect 31944 41550 31996 41556
rect 32220 41608 32272 41614
rect 32220 41550 32272 41556
rect 31850 41032 31906 41041
rect 31850 40967 31906 40976
rect 31760 40520 31812 40526
rect 31760 40462 31812 40468
rect 31576 40180 31628 40186
rect 31576 40122 31628 40128
rect 31588 38282 31616 40122
rect 31772 40118 31800 40462
rect 31864 40458 31892 40967
rect 31852 40452 31904 40458
rect 31852 40394 31904 40400
rect 31760 40112 31812 40118
rect 31760 40054 31812 40060
rect 31668 39092 31720 39098
rect 31668 39034 31720 39040
rect 31680 38282 31708 39034
rect 31772 38593 31800 40054
rect 31864 39642 31892 40394
rect 31852 39636 31904 39642
rect 31852 39578 31904 39584
rect 31758 38584 31814 38593
rect 31758 38519 31814 38528
rect 31852 38480 31904 38486
rect 31852 38422 31904 38428
rect 31576 38276 31628 38282
rect 31576 38218 31628 38224
rect 31668 38276 31720 38282
rect 31668 38218 31720 38224
rect 31484 38004 31536 38010
rect 31484 37946 31536 37952
rect 31392 36848 31444 36854
rect 31392 36790 31444 36796
rect 31496 36310 31524 37946
rect 31588 37874 31616 38218
rect 31576 37868 31628 37874
rect 31576 37810 31628 37816
rect 31484 36304 31536 36310
rect 31484 36246 31536 36252
rect 31392 36236 31444 36242
rect 31392 36178 31444 36184
rect 31300 35760 31352 35766
rect 31300 35702 31352 35708
rect 31208 35692 31260 35698
rect 31208 35634 31260 35640
rect 31220 35290 31248 35634
rect 31208 35284 31260 35290
rect 31208 35226 31260 35232
rect 31312 35086 31340 35702
rect 31404 35698 31432 36178
rect 31680 35834 31708 38218
rect 31864 38214 31892 38422
rect 31852 38208 31904 38214
rect 31852 38150 31904 38156
rect 31956 37942 31984 41550
rect 32312 41132 32364 41138
rect 32312 41074 32364 41080
rect 32324 39914 32352 41074
rect 32416 40730 32444 42026
rect 32404 40724 32456 40730
rect 32404 40666 32456 40672
rect 32416 40594 32444 40666
rect 32404 40588 32456 40594
rect 32404 40530 32456 40536
rect 32508 40050 32536 42638
rect 32692 42022 32720 42656
rect 32680 42016 32732 42022
rect 32680 41958 32732 41964
rect 32588 40452 32640 40458
rect 32692 40440 32720 41958
rect 32784 41614 32812 44814
rect 32876 44538 32904 44814
rect 32864 44532 32916 44538
rect 32864 44474 32916 44480
rect 32968 44334 32996 44934
rect 33060 44810 33088 45766
rect 33336 45490 33364 45970
rect 33416 45960 33468 45966
rect 33416 45902 33468 45908
rect 33428 45558 33456 45902
rect 33416 45552 33468 45558
rect 33416 45494 33468 45500
rect 33324 45484 33376 45490
rect 33324 45426 33376 45432
rect 33336 44860 33364 45426
rect 33508 44872 33560 44878
rect 33336 44832 33508 44860
rect 33048 44804 33100 44810
rect 33048 44746 33100 44752
rect 32956 44328 33008 44334
rect 32956 44270 33008 44276
rect 32956 43308 33008 43314
rect 32956 43250 33008 43256
rect 32864 43240 32916 43246
rect 32864 43182 32916 43188
rect 32772 41608 32824 41614
rect 32772 41550 32824 41556
rect 32784 41414 32812 41550
rect 32876 41546 32904 43182
rect 32968 42906 32996 43250
rect 32956 42900 33008 42906
rect 32956 42842 33008 42848
rect 33060 42634 33088 44746
rect 33336 44402 33364 44832
rect 33508 44814 33560 44820
rect 33324 44396 33376 44402
rect 33324 44338 33376 44344
rect 33336 43926 33364 44338
rect 33324 43920 33376 43926
rect 33324 43862 33376 43868
rect 33336 42906 33364 43862
rect 33612 43722 33640 46310
rect 33692 45892 33744 45898
rect 33692 45834 33744 45840
rect 33704 45626 33732 45834
rect 33796 45830 33824 46446
rect 34256 46034 34284 46582
rect 34244 46028 34296 46034
rect 34244 45970 34296 45976
rect 33784 45824 33836 45830
rect 33784 45766 33836 45772
rect 33692 45620 33744 45626
rect 33692 45562 33744 45568
rect 33796 44810 33824 45766
rect 34060 45076 34112 45082
rect 34060 45018 34112 45024
rect 33784 44804 33836 44810
rect 33784 44746 33836 44752
rect 33600 43716 33652 43722
rect 33600 43658 33652 43664
rect 33796 43654 33824 44746
rect 34072 44402 34100 45018
rect 34256 45014 34284 45970
rect 34336 45892 34388 45898
rect 34336 45834 34388 45840
rect 34348 45490 34376 45834
rect 34532 45626 34560 46854
rect 34716 46714 34744 48010
rect 34704 46708 34756 46714
rect 34704 46650 34756 46656
rect 34612 46572 34664 46578
rect 34612 46514 34664 46520
rect 34624 46170 34652 46514
rect 34612 46164 34664 46170
rect 34612 46106 34664 46112
rect 34808 45966 34836 48486
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 35072 48136 35124 48142
rect 35072 48078 35124 48084
rect 35084 47802 35112 48078
rect 35072 47796 35124 47802
rect 35072 47738 35124 47744
rect 35360 47530 35388 48690
rect 36268 48680 36320 48686
rect 36268 48622 36320 48628
rect 37556 48680 37608 48686
rect 37556 48622 37608 48628
rect 36280 48278 36308 48622
rect 37568 48278 37596 48622
rect 36268 48272 36320 48278
rect 36268 48214 36320 48220
rect 37556 48272 37608 48278
rect 37556 48214 37608 48220
rect 35992 48204 36044 48210
rect 35992 48146 36044 48152
rect 35594 47900 35902 47909
rect 35594 47898 35600 47900
rect 35656 47898 35680 47900
rect 35736 47898 35760 47900
rect 35816 47898 35840 47900
rect 35896 47898 35902 47900
rect 35656 47846 35658 47898
rect 35838 47846 35840 47898
rect 35594 47844 35600 47846
rect 35656 47844 35680 47846
rect 35736 47844 35760 47846
rect 35816 47844 35840 47846
rect 35896 47844 35902 47846
rect 35594 47835 35902 47844
rect 35624 47796 35676 47802
rect 35624 47738 35676 47744
rect 35532 47660 35584 47666
rect 35532 47602 35584 47608
rect 35348 47524 35400 47530
rect 35348 47466 35400 47472
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 35348 47048 35400 47054
rect 35348 46990 35400 46996
rect 35164 46980 35216 46986
rect 35164 46922 35216 46928
rect 35176 46646 35204 46922
rect 35164 46640 35216 46646
rect 35164 46582 35216 46588
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 35360 46102 35388 46990
rect 35544 46900 35572 47602
rect 35636 46918 35664 47738
rect 36004 47666 36032 48146
rect 36728 48068 36780 48074
rect 36728 48010 36780 48016
rect 36084 47728 36136 47734
rect 36084 47670 36136 47676
rect 35992 47660 36044 47666
rect 35992 47602 36044 47608
rect 35452 46872 35572 46900
rect 35624 46912 35676 46918
rect 35348 46096 35400 46102
rect 35348 46038 35400 46044
rect 34796 45960 34848 45966
rect 34796 45902 34848 45908
rect 34888 45960 34940 45966
rect 34888 45902 34940 45908
rect 34520 45620 34572 45626
rect 34520 45562 34572 45568
rect 34336 45484 34388 45490
rect 34336 45426 34388 45432
rect 34348 45014 34376 45426
rect 34520 45416 34572 45422
rect 34440 45364 34520 45370
rect 34440 45358 34572 45364
rect 34440 45342 34560 45358
rect 34900 45354 34928 45902
rect 35360 45830 35388 46038
rect 35348 45824 35400 45830
rect 35348 45766 35400 45772
rect 35452 45554 35480 46872
rect 35624 46854 35676 46860
rect 35594 46812 35902 46821
rect 35594 46810 35600 46812
rect 35656 46810 35680 46812
rect 35736 46810 35760 46812
rect 35816 46810 35840 46812
rect 35896 46810 35902 46812
rect 35656 46758 35658 46810
rect 35838 46758 35840 46810
rect 35594 46756 35600 46758
rect 35656 46756 35680 46758
rect 35736 46756 35760 46758
rect 35816 46756 35840 46758
rect 35896 46756 35902 46758
rect 35594 46747 35902 46756
rect 35532 46572 35584 46578
rect 35532 46514 35584 46520
rect 35544 46170 35572 46514
rect 35532 46164 35584 46170
rect 35532 46106 35584 46112
rect 35900 45960 35952 45966
rect 36004 45948 36032 47602
rect 36096 46578 36124 47670
rect 36740 47054 36768 48010
rect 36176 47048 36228 47054
rect 36176 46990 36228 46996
rect 36728 47048 36780 47054
rect 36728 46990 36780 46996
rect 37556 47048 37608 47054
rect 37556 46990 37608 46996
rect 36084 46572 36136 46578
rect 36084 46514 36136 46520
rect 35952 45920 36032 45948
rect 35900 45902 35952 45908
rect 35594 45724 35902 45733
rect 35594 45722 35600 45724
rect 35656 45722 35680 45724
rect 35736 45722 35760 45724
rect 35816 45722 35840 45724
rect 35896 45722 35902 45724
rect 35656 45670 35658 45722
rect 35838 45670 35840 45722
rect 35594 45668 35600 45670
rect 35656 45668 35680 45670
rect 35736 45668 35760 45670
rect 35816 45668 35840 45670
rect 35896 45668 35902 45670
rect 35594 45659 35902 45668
rect 35452 45526 35572 45554
rect 35440 45484 35492 45490
rect 35440 45426 35492 45432
rect 34888 45348 34940 45354
rect 34244 45008 34296 45014
rect 34244 44950 34296 44956
rect 34336 45008 34388 45014
rect 34336 44950 34388 44956
rect 34060 44396 34112 44402
rect 34060 44338 34112 44344
rect 34256 43994 34284 44950
rect 34440 44334 34468 45342
rect 34888 45290 34940 45296
rect 35348 45280 35400 45286
rect 35348 45222 35400 45228
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 35360 44946 35388 45222
rect 34612 44940 34664 44946
rect 34612 44882 34664 44888
rect 35348 44940 35400 44946
rect 35348 44882 35400 44888
rect 34520 44872 34572 44878
rect 34520 44814 34572 44820
rect 34532 44538 34560 44814
rect 34624 44742 34652 44882
rect 34612 44736 34664 44742
rect 34612 44678 34664 44684
rect 34520 44532 34572 44538
rect 34520 44474 34572 44480
rect 34520 44396 34572 44402
rect 34520 44338 34572 44344
rect 34428 44328 34480 44334
rect 34428 44270 34480 44276
rect 34244 43988 34296 43994
rect 34244 43930 34296 43936
rect 33784 43648 33836 43654
rect 33784 43590 33836 43596
rect 34060 43648 34112 43654
rect 34060 43590 34112 43596
rect 33968 43308 34020 43314
rect 33968 43250 34020 43256
rect 33980 43110 34008 43250
rect 34072 43246 34100 43590
rect 34060 43240 34112 43246
rect 34060 43182 34112 43188
rect 33968 43104 34020 43110
rect 33968 43046 34020 43052
rect 33324 42900 33376 42906
rect 33324 42842 33376 42848
rect 34072 42702 34100 43182
rect 34060 42696 34112 42702
rect 34060 42638 34112 42644
rect 33048 42628 33100 42634
rect 33048 42570 33100 42576
rect 32864 41540 32916 41546
rect 32864 41482 32916 41488
rect 32784 41386 32904 41414
rect 32772 40520 32824 40526
rect 32772 40462 32824 40468
rect 32640 40412 32720 40440
rect 32588 40394 32640 40400
rect 32496 40044 32548 40050
rect 32496 39986 32548 39992
rect 32312 39908 32364 39914
rect 32312 39850 32364 39856
rect 32220 39840 32272 39846
rect 32220 39782 32272 39788
rect 32232 39352 32260 39782
rect 32312 39364 32364 39370
rect 32232 39324 32312 39352
rect 32312 39306 32364 39312
rect 32324 38962 32352 39306
rect 32508 39098 32536 39986
rect 32600 39642 32628 40394
rect 32588 39636 32640 39642
rect 32588 39578 32640 39584
rect 32496 39092 32548 39098
rect 32496 39034 32548 39040
rect 32784 39030 32812 40462
rect 32772 39024 32824 39030
rect 32772 38966 32824 38972
rect 32312 38956 32364 38962
rect 32312 38898 32364 38904
rect 32680 38956 32732 38962
rect 32680 38898 32732 38904
rect 32220 38752 32272 38758
rect 32220 38694 32272 38700
rect 32232 38350 32260 38694
rect 32220 38344 32272 38350
rect 32220 38286 32272 38292
rect 31944 37936 31996 37942
rect 31944 37878 31996 37884
rect 32324 37466 32352 38898
rect 32692 38593 32720 38898
rect 32678 38584 32734 38593
rect 32678 38519 32734 38528
rect 32692 38350 32720 38519
rect 32496 38344 32548 38350
rect 32496 38286 32548 38292
rect 32680 38344 32732 38350
rect 32680 38286 32732 38292
rect 32508 37942 32536 38286
rect 32496 37936 32548 37942
rect 32496 37878 32548 37884
rect 32692 37466 32720 38286
rect 32784 37466 32812 38966
rect 32312 37460 32364 37466
rect 32312 37402 32364 37408
rect 32680 37460 32732 37466
rect 32680 37402 32732 37408
rect 32772 37460 32824 37466
rect 32772 37402 32824 37408
rect 32680 37324 32732 37330
rect 32876 37312 32904 41386
rect 32956 40384 33008 40390
rect 32956 40326 33008 40332
rect 32968 40050 32996 40326
rect 32956 40044 33008 40050
rect 32956 39986 33008 39992
rect 33060 38826 33088 42570
rect 34152 42220 34204 42226
rect 34152 42162 34204 42168
rect 33692 42084 33744 42090
rect 33692 42026 33744 42032
rect 33704 41818 33732 42026
rect 34164 42022 34192 42162
rect 34152 42016 34204 42022
rect 34150 41984 34152 41993
rect 34204 41984 34206 41993
rect 34150 41919 34206 41928
rect 33692 41812 33744 41818
rect 33692 41754 33744 41760
rect 33324 41676 33376 41682
rect 33324 41618 33376 41624
rect 33336 41138 33364 41618
rect 33968 41540 34020 41546
rect 33968 41482 34020 41488
rect 33324 41132 33376 41138
rect 33324 41074 33376 41080
rect 33232 40520 33284 40526
rect 33232 40462 33284 40468
rect 33244 40118 33272 40462
rect 33232 40112 33284 40118
rect 33232 40054 33284 40060
rect 33600 40044 33652 40050
rect 33600 39986 33652 39992
rect 33508 39976 33560 39982
rect 33508 39918 33560 39924
rect 33520 39438 33548 39918
rect 33508 39432 33560 39438
rect 33508 39374 33560 39380
rect 33612 38962 33640 39986
rect 33980 39914 34008 41482
rect 34256 41414 34284 43930
rect 34440 43858 34468 44270
rect 34428 43852 34480 43858
rect 34428 43794 34480 43800
rect 34336 43716 34388 43722
rect 34336 43658 34388 43664
rect 34164 41386 34284 41414
rect 34060 39976 34112 39982
rect 34060 39918 34112 39924
rect 33968 39908 34020 39914
rect 33968 39850 34020 39856
rect 34072 39642 34100 39918
rect 34060 39636 34112 39642
rect 34060 39578 34112 39584
rect 33876 39500 33928 39506
rect 33876 39442 33928 39448
rect 33600 38956 33652 38962
rect 33600 38898 33652 38904
rect 33048 38820 33100 38826
rect 33048 38762 33100 38768
rect 33060 38010 33088 38762
rect 33416 38412 33468 38418
rect 33416 38354 33468 38360
rect 33048 38004 33100 38010
rect 33048 37946 33100 37952
rect 32876 37284 33088 37312
rect 32680 37266 32732 37272
rect 32692 36786 32720 37266
rect 32956 37188 33008 37194
rect 32956 37130 33008 37136
rect 32968 36854 32996 37130
rect 32864 36848 32916 36854
rect 32864 36790 32916 36796
rect 32956 36848 33008 36854
rect 32956 36790 33008 36796
rect 32680 36780 32732 36786
rect 32680 36722 32732 36728
rect 32772 36780 32824 36786
rect 32772 36722 32824 36728
rect 32496 36032 32548 36038
rect 32496 35974 32548 35980
rect 31668 35828 31720 35834
rect 31668 35770 31720 35776
rect 31392 35692 31444 35698
rect 31392 35634 31444 35640
rect 31680 35170 31708 35770
rect 32312 35488 32364 35494
rect 32312 35430 32364 35436
rect 32404 35488 32456 35494
rect 32404 35430 32456 35436
rect 32036 35284 32088 35290
rect 32036 35226 32088 35232
rect 31680 35142 31984 35170
rect 31300 35080 31352 35086
rect 31300 35022 31352 35028
rect 31760 35080 31812 35086
rect 31760 35022 31812 35028
rect 31208 35012 31260 35018
rect 31208 34954 31260 34960
rect 31220 34610 31248 34954
rect 31772 34678 31800 35022
rect 31956 34678 31984 35142
rect 32048 35018 32076 35226
rect 32036 35012 32088 35018
rect 32036 34954 32088 34960
rect 31760 34672 31812 34678
rect 31760 34614 31812 34620
rect 31944 34672 31996 34678
rect 31944 34614 31996 34620
rect 31208 34604 31260 34610
rect 31208 34546 31260 34552
rect 30288 32020 30340 32026
rect 30288 31962 30340 31968
rect 31116 32020 31168 32026
rect 31116 31962 31168 31968
rect 30196 31952 30248 31958
rect 30196 31894 30248 31900
rect 29828 31680 29880 31686
rect 29828 31622 29880 31628
rect 29840 31414 29868 31622
rect 29828 31408 29880 31414
rect 29828 31350 29880 31356
rect 30208 31346 30236 31894
rect 30300 31822 30328 31962
rect 30288 31816 30340 31822
rect 30288 31758 30340 31764
rect 30196 31340 30248 31346
rect 30196 31282 30248 31288
rect 29460 30796 29512 30802
rect 29460 30738 29512 30744
rect 30300 30258 30328 31758
rect 30840 30660 30892 30666
rect 30840 30602 30892 30608
rect 30852 30326 30880 30602
rect 30840 30320 30892 30326
rect 30840 30262 30892 30268
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 29368 29844 29420 29850
rect 29368 29786 29420 29792
rect 30196 29640 30248 29646
rect 30196 29582 30248 29588
rect 28816 29504 28868 29510
rect 28816 29446 28868 29452
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 30208 29306 30236 29582
rect 30196 29300 30248 29306
rect 30196 29242 30248 29248
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 31220 28762 31248 34546
rect 31668 34536 31720 34542
rect 31668 34478 31720 34484
rect 31680 33998 31708 34478
rect 31668 33992 31720 33998
rect 31668 33934 31720 33940
rect 31772 33590 31800 34614
rect 32324 34406 32352 35430
rect 32416 35086 32444 35430
rect 32404 35080 32456 35086
rect 32404 35022 32456 35028
rect 32508 34746 32536 35974
rect 32784 35562 32812 36722
rect 32876 35630 32904 36790
rect 33060 36242 33088 37284
rect 33140 37188 33192 37194
rect 33140 37130 33192 37136
rect 33152 36582 33180 37130
rect 33140 36576 33192 36582
rect 33140 36518 33192 36524
rect 33152 36378 33180 36518
rect 33140 36372 33192 36378
rect 33140 36314 33192 36320
rect 33048 36236 33100 36242
rect 33048 36178 33100 36184
rect 33322 36136 33378 36145
rect 33322 36071 33324 36080
rect 33376 36071 33378 36080
rect 33324 36042 33376 36048
rect 33324 35692 33376 35698
rect 33324 35634 33376 35640
rect 32864 35624 32916 35630
rect 32864 35566 32916 35572
rect 32772 35556 32824 35562
rect 32772 35498 32824 35504
rect 32956 35556 33008 35562
rect 32956 35498 33008 35504
rect 32784 35222 32812 35498
rect 32772 35216 32824 35222
rect 32772 35158 32824 35164
rect 32772 35080 32824 35086
rect 32968 35034 32996 35498
rect 33336 35086 33364 35634
rect 32824 35028 32996 35034
rect 32772 35022 32996 35028
rect 33324 35080 33376 35086
rect 33324 35022 33376 35028
rect 32784 35006 32996 35022
rect 32680 34944 32732 34950
rect 32680 34886 32732 34892
rect 32692 34746 32720 34886
rect 32496 34740 32548 34746
rect 32496 34682 32548 34688
rect 32680 34740 32732 34746
rect 32680 34682 32732 34688
rect 32784 34406 32812 35006
rect 33232 34672 33284 34678
rect 33232 34614 33284 34620
rect 33140 34604 33192 34610
rect 33140 34546 33192 34552
rect 32312 34400 32364 34406
rect 32312 34342 32364 34348
rect 32772 34400 32824 34406
rect 32772 34342 32824 34348
rect 33048 34400 33100 34406
rect 33048 34342 33100 34348
rect 33060 33998 33088 34342
rect 33152 34202 33180 34546
rect 33140 34196 33192 34202
rect 33140 34138 33192 34144
rect 33048 33992 33100 33998
rect 33048 33934 33100 33940
rect 31760 33584 31812 33590
rect 31760 33526 31812 33532
rect 33060 33454 33088 33934
rect 33244 33522 33272 34614
rect 33336 33930 33364 35022
rect 33428 34474 33456 38354
rect 33508 37936 33560 37942
rect 33508 37878 33560 37884
rect 33520 37262 33548 37878
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 33508 36168 33560 36174
rect 33508 36110 33560 36116
rect 33520 35290 33548 36110
rect 33612 35766 33640 38898
rect 33888 38894 33916 39442
rect 33876 38888 33928 38894
rect 33690 38856 33746 38865
rect 33876 38830 33928 38836
rect 33690 38791 33746 38800
rect 33704 38418 33732 38791
rect 33888 38554 33916 38830
rect 33876 38548 33928 38554
rect 33876 38490 33928 38496
rect 33692 38412 33744 38418
rect 33692 38354 33744 38360
rect 33692 37936 33744 37942
rect 33692 37878 33744 37884
rect 33704 37262 33732 37878
rect 33784 37664 33836 37670
rect 33784 37606 33836 37612
rect 33692 37256 33744 37262
rect 33692 37198 33744 37204
rect 33704 36689 33732 37198
rect 33796 37194 33824 37606
rect 34164 37482 34192 41386
rect 34072 37454 34192 37482
rect 34072 37398 34100 37454
rect 34060 37392 34112 37398
rect 34060 37334 34112 37340
rect 33876 37324 33928 37330
rect 33876 37266 33928 37272
rect 33888 37194 33916 37266
rect 33784 37188 33836 37194
rect 33784 37130 33836 37136
rect 33876 37188 33928 37194
rect 33876 37130 33928 37136
rect 33796 36922 33824 37130
rect 33784 36916 33836 36922
rect 33784 36858 33836 36864
rect 33690 36680 33746 36689
rect 34072 36666 34100 37334
rect 34348 37312 34376 43658
rect 34532 43450 34560 44338
rect 34520 43444 34572 43450
rect 34520 43386 34572 43392
rect 34624 42226 34652 44678
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 35348 43920 35400 43926
rect 35348 43862 35400 43868
rect 35072 43716 35124 43722
rect 35072 43658 35124 43664
rect 35084 43314 35112 43658
rect 35360 43450 35388 43862
rect 35348 43444 35400 43450
rect 35348 43386 35400 43392
rect 34796 43308 34848 43314
rect 34796 43250 34848 43256
rect 35072 43308 35124 43314
rect 35072 43250 35124 43256
rect 35256 43308 35308 43314
rect 35308 43268 35388 43296
rect 35256 43250 35308 43256
rect 34704 42832 34756 42838
rect 34704 42774 34756 42780
rect 34716 42226 34744 42774
rect 34808 42362 34836 43250
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34980 42764 35032 42770
rect 34980 42706 35032 42712
rect 34888 42560 34940 42566
rect 34888 42502 34940 42508
rect 34796 42356 34848 42362
rect 34796 42298 34848 42304
rect 34900 42242 34928 42502
rect 34992 42362 35020 42706
rect 35256 42696 35308 42702
rect 35256 42638 35308 42644
rect 35268 42514 35296 42638
rect 35360 42634 35388 43268
rect 35348 42628 35400 42634
rect 35348 42570 35400 42576
rect 35452 42548 35480 45426
rect 35544 44878 35572 45526
rect 36188 45354 36216 46990
rect 36452 46436 36504 46442
rect 36452 46378 36504 46384
rect 36464 46034 36492 46378
rect 36452 46028 36504 46034
rect 36452 45970 36504 45976
rect 36740 45966 36768 46990
rect 37464 46980 37516 46986
rect 37464 46922 37516 46928
rect 37476 46578 37504 46922
rect 37568 46594 37596 46990
rect 37660 46714 37688 48690
rect 38752 48680 38804 48686
rect 38752 48622 38804 48628
rect 38476 48612 38528 48618
rect 38476 48554 38528 48560
rect 38488 48278 38516 48554
rect 38764 48550 38792 48622
rect 38752 48544 38804 48550
rect 38752 48486 38804 48492
rect 38476 48272 38528 48278
rect 38476 48214 38528 48220
rect 38764 48142 38792 48486
rect 40132 48204 40184 48210
rect 40132 48146 40184 48152
rect 38752 48136 38804 48142
rect 38752 48078 38804 48084
rect 38292 48000 38344 48006
rect 38292 47942 38344 47948
rect 37740 47592 37792 47598
rect 37740 47534 37792 47540
rect 37648 46708 37700 46714
rect 37648 46650 37700 46656
rect 37568 46578 37688 46594
rect 37464 46572 37516 46578
rect 37568 46572 37700 46578
rect 37568 46566 37648 46572
rect 37464 46514 37516 46520
rect 37648 46514 37700 46520
rect 37372 46436 37424 46442
rect 37372 46378 37424 46384
rect 36360 45960 36412 45966
rect 36360 45902 36412 45908
rect 36728 45960 36780 45966
rect 36728 45902 36780 45908
rect 36372 45626 36400 45902
rect 36360 45620 36412 45626
rect 36360 45562 36412 45568
rect 36176 45348 36228 45354
rect 36176 45290 36228 45296
rect 36188 45098 36216 45290
rect 36096 45070 36216 45098
rect 36096 45014 36124 45070
rect 36084 45008 36136 45014
rect 36084 44950 36136 44956
rect 35532 44872 35584 44878
rect 35532 44814 35584 44820
rect 35594 44636 35902 44645
rect 35594 44634 35600 44636
rect 35656 44634 35680 44636
rect 35736 44634 35760 44636
rect 35816 44634 35840 44636
rect 35896 44634 35902 44636
rect 35656 44582 35658 44634
rect 35838 44582 35840 44634
rect 35594 44580 35600 44582
rect 35656 44580 35680 44582
rect 35736 44580 35760 44582
rect 35816 44580 35840 44582
rect 35896 44580 35902 44582
rect 35594 44571 35902 44580
rect 36372 43994 36400 45562
rect 36636 45484 36688 45490
rect 36636 45426 36688 45432
rect 36648 44402 36676 45426
rect 36912 44872 36964 44878
rect 36912 44814 36964 44820
rect 36636 44396 36688 44402
rect 36636 44338 36688 44344
rect 36924 44266 36952 44814
rect 37188 44328 37240 44334
rect 37240 44288 37320 44316
rect 37188 44270 37240 44276
rect 36912 44260 36964 44266
rect 36912 44202 36964 44208
rect 36728 44192 36780 44198
rect 36728 44134 36780 44140
rect 36360 43988 36412 43994
rect 36412 43948 36492 43976
rect 36360 43930 36412 43936
rect 36268 43920 36320 43926
rect 36268 43862 36320 43868
rect 35594 43548 35902 43557
rect 35594 43546 35600 43548
rect 35656 43546 35680 43548
rect 35736 43546 35760 43548
rect 35816 43546 35840 43548
rect 35896 43546 35902 43548
rect 35656 43494 35658 43546
rect 35838 43494 35840 43546
rect 35594 43492 35600 43494
rect 35656 43492 35680 43494
rect 35736 43492 35760 43494
rect 35816 43492 35840 43494
rect 35896 43492 35902 43494
rect 35594 43483 35902 43492
rect 36084 43444 36136 43450
rect 36084 43386 36136 43392
rect 36096 43353 36124 43386
rect 36176 43376 36228 43382
rect 36082 43344 36138 43353
rect 35532 43308 35584 43314
rect 36176 43318 36228 43324
rect 36082 43279 36138 43288
rect 35532 43250 35584 43256
rect 35544 42702 35572 43250
rect 35624 43240 35676 43246
rect 35624 43182 35676 43188
rect 35532 42696 35584 42702
rect 35532 42638 35584 42644
rect 35636 42634 35664 43182
rect 35992 42696 36044 42702
rect 35992 42638 36044 42644
rect 35624 42628 35676 42634
rect 35624 42570 35676 42576
rect 35532 42560 35584 42566
rect 35452 42520 35532 42548
rect 35268 42486 35388 42514
rect 35532 42502 35584 42508
rect 35360 42378 35388 42486
rect 35594 42460 35902 42469
rect 35594 42458 35600 42460
rect 35656 42458 35680 42460
rect 35736 42458 35760 42460
rect 35816 42458 35840 42460
rect 35896 42458 35902 42460
rect 35656 42406 35658 42458
rect 35838 42406 35840 42458
rect 35594 42404 35600 42406
rect 35656 42404 35680 42406
rect 35736 42404 35760 42406
rect 35816 42404 35840 42406
rect 35896 42404 35902 42406
rect 35594 42395 35902 42404
rect 34980 42356 35032 42362
rect 35360 42350 35480 42378
rect 36004 42362 36032 42638
rect 34980 42298 35032 42304
rect 34612 42220 34664 42226
rect 34612 42162 34664 42168
rect 34704 42220 34756 42226
rect 34704 42162 34756 42168
rect 34808 42214 34928 42242
rect 34716 41682 34744 42162
rect 34704 41676 34756 41682
rect 34704 41618 34756 41624
rect 34716 40730 34744 41618
rect 34808 41206 34836 42214
rect 34992 42158 35020 42298
rect 35452 42158 35480 42350
rect 35992 42356 36044 42362
rect 35992 42298 36044 42304
rect 36096 42226 36124 43279
rect 36188 42566 36216 43318
rect 36176 42560 36228 42566
rect 36176 42502 36228 42508
rect 36188 42294 36216 42502
rect 36176 42288 36228 42294
rect 36176 42230 36228 42236
rect 36084 42220 36136 42226
rect 36084 42162 36136 42168
rect 34980 42152 35032 42158
rect 34980 42094 35032 42100
rect 35348 42152 35400 42158
rect 35348 42094 35400 42100
rect 35440 42152 35492 42158
rect 35440 42094 35492 42100
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34980 41608 35032 41614
rect 34980 41550 35032 41556
rect 34992 41274 35020 41550
rect 34980 41268 35032 41274
rect 34980 41210 35032 41216
rect 34796 41200 34848 41206
rect 34796 41142 34848 41148
rect 34704 40724 34756 40730
rect 34704 40666 34756 40672
rect 34612 40112 34664 40118
rect 34612 40054 34664 40060
rect 34428 39296 34480 39302
rect 34428 39238 34480 39244
rect 34440 39098 34468 39238
rect 34428 39092 34480 39098
rect 34428 39034 34480 39040
rect 34624 38962 34652 40054
rect 34612 38956 34664 38962
rect 34612 38898 34664 38904
rect 34624 38486 34652 38898
rect 34716 38894 34744 40666
rect 34808 39370 34836 41142
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35360 40594 35388 42094
rect 35452 41138 35480 42094
rect 35594 41372 35902 41381
rect 35594 41370 35600 41372
rect 35656 41370 35680 41372
rect 35736 41370 35760 41372
rect 35816 41370 35840 41372
rect 35896 41370 35902 41372
rect 35656 41318 35658 41370
rect 35838 41318 35840 41370
rect 35594 41316 35600 41318
rect 35656 41316 35680 41318
rect 35736 41316 35760 41318
rect 35816 41316 35840 41318
rect 35896 41316 35902 41318
rect 35594 41307 35902 41316
rect 35440 41132 35492 41138
rect 35440 41074 35492 41080
rect 35532 41132 35584 41138
rect 35532 41074 35584 41080
rect 35808 41132 35860 41138
rect 35808 41074 35860 41080
rect 35900 41132 35952 41138
rect 35900 41074 35952 41080
rect 35452 41002 35480 41074
rect 35440 40996 35492 41002
rect 35440 40938 35492 40944
rect 35544 40662 35572 41074
rect 35820 41041 35848 41074
rect 35806 41032 35862 41041
rect 35806 40967 35862 40976
rect 35912 40730 35940 41074
rect 35992 40996 36044 41002
rect 35992 40938 36044 40944
rect 35900 40724 35952 40730
rect 35900 40666 35952 40672
rect 35532 40656 35584 40662
rect 35532 40598 35584 40604
rect 35348 40588 35400 40594
rect 35348 40530 35400 40536
rect 35256 40520 35308 40526
rect 35256 40462 35308 40468
rect 35268 39846 35296 40462
rect 35256 39840 35308 39846
rect 35256 39782 35308 39788
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 35256 39500 35308 39506
rect 35256 39442 35308 39448
rect 34796 39364 34848 39370
rect 34796 39306 34848 39312
rect 34704 38888 34756 38894
rect 34704 38830 34756 38836
rect 34612 38480 34664 38486
rect 34612 38422 34664 38428
rect 34520 38344 34572 38350
rect 34520 38286 34572 38292
rect 33690 36615 33746 36624
rect 33888 36638 34100 36666
rect 34164 37284 34376 37312
rect 33692 36304 33744 36310
rect 33692 36246 33744 36252
rect 33600 35760 33652 35766
rect 33600 35702 33652 35708
rect 33508 35284 33560 35290
rect 33508 35226 33560 35232
rect 33704 35086 33732 36246
rect 33888 36122 33916 36638
rect 33968 36576 34020 36582
rect 33968 36518 34020 36524
rect 33796 36106 33916 36122
rect 33784 36100 33916 36106
rect 33836 36094 33916 36100
rect 33784 36042 33836 36048
rect 33782 36000 33838 36009
rect 33782 35935 33838 35944
rect 33692 35080 33744 35086
rect 33692 35022 33744 35028
rect 33796 35018 33824 35935
rect 33888 35290 33916 36094
rect 33876 35284 33928 35290
rect 33876 35226 33928 35232
rect 33980 35222 34008 36518
rect 34060 36372 34112 36378
rect 34060 36314 34112 36320
rect 34072 36242 34100 36314
rect 34060 36236 34112 36242
rect 34060 36178 34112 36184
rect 34060 36032 34112 36038
rect 34060 35974 34112 35980
rect 34072 35698 34100 35974
rect 34060 35692 34112 35698
rect 34060 35634 34112 35640
rect 33968 35216 34020 35222
rect 33968 35158 34020 35164
rect 33784 35012 33836 35018
rect 33784 34954 33836 34960
rect 33796 34610 33824 34954
rect 33784 34604 33836 34610
rect 33784 34546 33836 34552
rect 33416 34468 33468 34474
rect 33416 34410 33468 34416
rect 33600 33992 33652 33998
rect 33600 33934 33652 33940
rect 33784 33992 33836 33998
rect 33784 33934 33836 33940
rect 33324 33924 33376 33930
rect 33324 33866 33376 33872
rect 33612 33658 33640 33934
rect 33600 33652 33652 33658
rect 33600 33594 33652 33600
rect 33796 33590 33824 33934
rect 33784 33584 33836 33590
rect 33784 33526 33836 33532
rect 33232 33516 33284 33522
rect 33232 33458 33284 33464
rect 33048 33448 33100 33454
rect 33048 33390 33100 33396
rect 34164 33114 34192 37284
rect 34428 37120 34480 37126
rect 34428 37062 34480 37068
rect 34440 36786 34468 37062
rect 34428 36780 34480 36786
rect 34428 36722 34480 36728
rect 34244 36712 34296 36718
rect 34244 36654 34296 36660
rect 34256 36378 34284 36654
rect 34244 36372 34296 36378
rect 34244 36314 34296 36320
rect 34532 34950 34560 38286
rect 34808 38010 34836 39306
rect 35268 38962 35296 39442
rect 35360 38978 35388 40530
rect 35594 40284 35902 40293
rect 35594 40282 35600 40284
rect 35656 40282 35680 40284
rect 35736 40282 35760 40284
rect 35816 40282 35840 40284
rect 35896 40282 35902 40284
rect 35656 40230 35658 40282
rect 35838 40230 35840 40282
rect 35594 40228 35600 40230
rect 35656 40228 35680 40230
rect 35736 40228 35760 40230
rect 35816 40228 35840 40230
rect 35896 40228 35902 40230
rect 35594 40219 35902 40228
rect 35532 39840 35584 39846
rect 35532 39782 35584 39788
rect 35544 39438 35572 39782
rect 36004 39438 36032 40938
rect 36084 40044 36136 40050
rect 36084 39986 36136 39992
rect 36096 39642 36124 39986
rect 36084 39636 36136 39642
rect 36084 39578 36136 39584
rect 35440 39432 35492 39438
rect 35440 39374 35492 39380
rect 35532 39432 35584 39438
rect 35532 39374 35584 39380
rect 35992 39432 36044 39438
rect 35992 39374 36044 39380
rect 35452 39098 35480 39374
rect 35594 39196 35902 39205
rect 35594 39194 35600 39196
rect 35656 39194 35680 39196
rect 35736 39194 35760 39196
rect 35816 39194 35840 39196
rect 35896 39194 35902 39196
rect 35656 39142 35658 39194
rect 35838 39142 35840 39194
rect 35594 39140 35600 39142
rect 35656 39140 35680 39142
rect 35736 39140 35760 39142
rect 35816 39140 35840 39142
rect 35896 39140 35902 39142
rect 35594 39131 35902 39140
rect 35440 39092 35492 39098
rect 35440 39034 35492 39040
rect 35256 38956 35308 38962
rect 35360 38950 35480 38978
rect 35256 38898 35308 38904
rect 35452 38894 35480 38950
rect 35348 38888 35400 38894
rect 35348 38830 35400 38836
rect 35440 38888 35492 38894
rect 35440 38830 35492 38836
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 35360 38554 35388 38830
rect 35452 38554 35480 38830
rect 35348 38548 35400 38554
rect 35348 38490 35400 38496
rect 35440 38548 35492 38554
rect 35440 38490 35492 38496
rect 35072 38344 35124 38350
rect 35072 38286 35124 38292
rect 34980 38276 35032 38282
rect 34980 38218 35032 38224
rect 34796 38004 34848 38010
rect 34796 37946 34848 37952
rect 34992 37874 35020 38218
rect 35084 38214 35112 38286
rect 35072 38208 35124 38214
rect 35072 38150 35124 38156
rect 35594 38108 35902 38117
rect 35594 38106 35600 38108
rect 35656 38106 35680 38108
rect 35736 38106 35760 38108
rect 35816 38106 35840 38108
rect 35896 38106 35902 38108
rect 35656 38054 35658 38106
rect 35838 38054 35840 38106
rect 35594 38052 35600 38054
rect 35656 38052 35680 38054
rect 35736 38052 35760 38054
rect 35816 38052 35840 38054
rect 35896 38052 35902 38054
rect 35594 38043 35902 38052
rect 36004 37942 36032 39374
rect 35532 37936 35584 37942
rect 35532 37878 35584 37884
rect 35992 37936 36044 37942
rect 35992 37878 36044 37884
rect 34980 37868 35032 37874
rect 34808 37828 34980 37856
rect 34612 37256 34664 37262
rect 34612 37198 34664 37204
rect 34624 36786 34652 37198
rect 34612 36780 34664 36786
rect 34612 36722 34664 36728
rect 34624 36038 34652 36722
rect 34612 36032 34664 36038
rect 34612 35974 34664 35980
rect 34520 34944 34572 34950
rect 34520 34886 34572 34892
rect 34336 34536 34388 34542
rect 34336 34478 34388 34484
rect 34348 34066 34376 34478
rect 34336 34060 34388 34066
rect 34336 34002 34388 34008
rect 34152 33108 34204 33114
rect 34152 33050 34204 33056
rect 32864 32904 32916 32910
rect 32864 32846 32916 32852
rect 31576 32836 31628 32842
rect 31576 32778 31628 32784
rect 31588 32570 31616 32778
rect 32876 32570 32904 32846
rect 31576 32564 31628 32570
rect 31576 32506 31628 32512
rect 32864 32564 32916 32570
rect 32864 32506 32916 32512
rect 32312 32360 32364 32366
rect 32312 32302 32364 32308
rect 32324 32026 32352 32302
rect 32312 32020 32364 32026
rect 32312 31962 32364 31968
rect 32404 31748 32456 31754
rect 32404 31690 32456 31696
rect 32680 31748 32732 31754
rect 32680 31690 32732 31696
rect 32416 31482 32444 31690
rect 32692 31482 32720 31690
rect 32404 31476 32456 31482
rect 32404 31418 32456 31424
rect 32680 31476 32732 31482
rect 32680 31418 32732 31424
rect 32876 31346 32904 32506
rect 34244 32496 34296 32502
rect 34244 32438 34296 32444
rect 32956 32360 33008 32366
rect 32956 32302 33008 32308
rect 32968 31890 32996 32302
rect 34256 32026 34284 32438
rect 34244 32020 34296 32026
rect 34244 31962 34296 31968
rect 32956 31884 33008 31890
rect 32956 31826 33008 31832
rect 32968 31346 32996 31826
rect 33876 31408 33928 31414
rect 33876 31350 33928 31356
rect 32864 31340 32916 31346
rect 32864 31282 32916 31288
rect 32956 31340 33008 31346
rect 32956 31282 33008 31288
rect 31852 30728 31904 30734
rect 31852 30670 31904 30676
rect 31668 30660 31720 30666
rect 31668 30602 31720 30608
rect 31680 29646 31708 30602
rect 31760 30252 31812 30258
rect 31760 30194 31812 30200
rect 31772 30054 31800 30194
rect 31760 30048 31812 30054
rect 31760 29990 31812 29996
rect 31668 29640 31720 29646
rect 31668 29582 31720 29588
rect 31300 29572 31352 29578
rect 31300 29514 31352 29520
rect 31312 29209 31340 29514
rect 31298 29200 31354 29209
rect 31772 29170 31800 29990
rect 31864 29850 31892 30670
rect 32402 30288 32458 30297
rect 32402 30223 32458 30232
rect 32772 30252 32824 30258
rect 32416 30054 32444 30223
rect 32772 30194 32824 30200
rect 32404 30048 32456 30054
rect 32404 29990 32456 29996
rect 31852 29844 31904 29850
rect 31852 29786 31904 29792
rect 32784 29306 32812 30194
rect 32772 29300 32824 29306
rect 32772 29242 32824 29248
rect 32876 29170 32904 31282
rect 33692 31272 33744 31278
rect 33692 31214 33744 31220
rect 33704 30938 33732 31214
rect 33692 30932 33744 30938
rect 33692 30874 33744 30880
rect 33888 30870 33916 31350
rect 33968 31136 34020 31142
rect 33968 31078 34020 31084
rect 33876 30864 33928 30870
rect 33876 30806 33928 30812
rect 33980 30734 34008 31078
rect 34348 30841 34376 34002
rect 34334 30832 34390 30841
rect 34334 30767 34390 30776
rect 33968 30728 34020 30734
rect 33968 30670 34020 30676
rect 34152 30728 34204 30734
rect 34152 30670 34204 30676
rect 34164 30258 34192 30670
rect 34152 30252 34204 30258
rect 34152 30194 34204 30200
rect 34164 29850 34192 30194
rect 34532 30138 34560 34886
rect 34624 33318 34652 35974
rect 34704 35828 34756 35834
rect 34704 35770 34756 35776
rect 34716 33658 34744 35770
rect 34704 33652 34756 33658
rect 34704 33594 34756 33600
rect 34704 33516 34756 33522
rect 34704 33458 34756 33464
rect 34612 33312 34664 33318
rect 34612 33254 34664 33260
rect 34624 33114 34652 33254
rect 34612 33108 34664 33114
rect 34612 33050 34664 33056
rect 34716 32570 34744 33458
rect 34808 32994 34836 37828
rect 35440 37868 35492 37874
rect 34980 37810 35032 37816
rect 35360 37828 35440 37856
rect 35360 37670 35388 37828
rect 35440 37810 35492 37816
rect 35348 37664 35400 37670
rect 35348 37606 35400 37612
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34888 36100 34940 36106
rect 34888 36042 34940 36048
rect 34900 35766 34928 36042
rect 34888 35760 34940 35766
rect 34888 35702 34940 35708
rect 35360 35630 35388 37606
rect 35544 37108 35572 37878
rect 35624 37392 35676 37398
rect 35624 37334 35676 37340
rect 35636 37126 35664 37334
rect 35992 37256 36044 37262
rect 35992 37198 36044 37204
rect 35452 37080 35572 37108
rect 35624 37120 35676 37126
rect 35452 35680 35480 37080
rect 35624 37062 35676 37068
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 35808 36916 35860 36922
rect 35808 36858 35860 36864
rect 35820 36718 35848 36858
rect 36004 36786 36032 37198
rect 35992 36780 36044 36786
rect 35992 36722 36044 36728
rect 35808 36712 35860 36718
rect 35808 36654 35860 36660
rect 35898 36680 35954 36689
rect 35898 36615 35954 36624
rect 35912 36038 35940 36615
rect 36004 36174 36032 36722
rect 36176 36644 36228 36650
rect 36176 36586 36228 36592
rect 35992 36168 36044 36174
rect 36044 36128 36124 36156
rect 35992 36110 36044 36116
rect 35900 36032 35952 36038
rect 35952 35992 36032 36020
rect 35900 35974 35952 35980
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 35716 35828 35768 35834
rect 36004 35816 36032 35992
rect 35768 35788 36032 35816
rect 35716 35770 35768 35776
rect 35452 35652 35848 35680
rect 35348 35624 35400 35630
rect 35348 35566 35400 35572
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35360 34678 35388 35566
rect 35440 35556 35492 35562
rect 35440 35498 35492 35504
rect 35452 35290 35480 35498
rect 35440 35284 35492 35290
rect 35440 35226 35492 35232
rect 35716 35080 35768 35086
rect 35452 35028 35716 35034
rect 35452 35022 35768 35028
rect 35452 35006 35756 35022
rect 35452 34950 35480 35006
rect 35820 34950 35848 35652
rect 35440 34944 35492 34950
rect 35440 34886 35492 34892
rect 35808 34944 35860 34950
rect 35860 34904 36032 34932
rect 35808 34886 35860 34892
rect 35348 34672 35400 34678
rect 35348 34614 35400 34620
rect 35452 34626 35480 34886
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 35452 34610 35572 34626
rect 35452 34604 35584 34610
rect 35452 34598 35532 34604
rect 35532 34546 35584 34552
rect 35348 34536 35400 34542
rect 35348 34478 35400 34484
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35360 33114 35388 34478
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 35440 33380 35492 33386
rect 35440 33322 35492 33328
rect 35348 33108 35400 33114
rect 35348 33050 35400 33056
rect 34808 32966 34928 32994
rect 34796 32904 34848 32910
rect 34796 32846 34848 32852
rect 34704 32564 34756 32570
rect 34704 32506 34756 32512
rect 34612 31884 34664 31890
rect 34612 31826 34664 31832
rect 34624 31414 34652 31826
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 34612 31408 34664 31414
rect 34612 31350 34664 31356
rect 34716 30682 34744 31758
rect 34808 30802 34836 32846
rect 34900 32434 34928 32966
rect 34888 32428 34940 32434
rect 34888 32370 34940 32376
rect 35348 32224 35400 32230
rect 35348 32166 35400 32172
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35360 32026 35388 32166
rect 35348 32020 35400 32026
rect 35348 31962 35400 31968
rect 35348 31884 35400 31890
rect 35348 31826 35400 31832
rect 35360 31482 35388 31826
rect 35348 31476 35400 31482
rect 35348 31418 35400 31424
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34796 30796 34848 30802
rect 34796 30738 34848 30744
rect 35348 30796 35400 30802
rect 35348 30738 35400 30744
rect 34716 30654 35020 30682
rect 34796 30592 34848 30598
rect 34796 30534 34848 30540
rect 34808 30394 34836 30534
rect 34704 30388 34756 30394
rect 34704 30330 34756 30336
rect 34796 30388 34848 30394
rect 34796 30330 34848 30336
rect 34716 30274 34744 30330
rect 34716 30246 34928 30274
rect 34900 30190 34928 30246
rect 34888 30184 34940 30190
rect 34532 30110 34652 30138
rect 34888 30126 34940 30132
rect 34520 30048 34572 30054
rect 34520 29990 34572 29996
rect 33416 29844 33468 29850
rect 33416 29786 33468 29792
rect 34152 29844 34204 29850
rect 34152 29786 34204 29792
rect 32956 29572 33008 29578
rect 32956 29514 33008 29520
rect 31298 29135 31354 29144
rect 31760 29164 31812 29170
rect 31760 29106 31812 29112
rect 32864 29164 32916 29170
rect 32864 29106 32916 29112
rect 31668 28960 31720 28966
rect 31668 28902 31720 28908
rect 31208 28756 31260 28762
rect 31208 28698 31260 28704
rect 31680 28490 31708 28902
rect 31668 28484 31720 28490
rect 31668 28426 31720 28432
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 31772 27878 31800 29106
rect 32312 28620 32364 28626
rect 32312 28562 32364 28568
rect 32324 28014 32352 28562
rect 32876 28558 32904 29106
rect 32864 28552 32916 28558
rect 32864 28494 32916 28500
rect 32312 28008 32364 28014
rect 32312 27950 32364 27956
rect 32588 28008 32640 28014
rect 32588 27950 32640 27956
rect 31760 27872 31812 27878
rect 31760 27814 31812 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 2412 26580 2464 26586
rect 2412 26522 2464 26528
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 31772 25294 31800 27814
rect 32324 26586 32352 27950
rect 32600 27674 32628 27950
rect 32968 27878 32996 29514
rect 33428 29170 33456 29786
rect 34336 29572 34388 29578
rect 34336 29514 34388 29520
rect 33416 29164 33468 29170
rect 33416 29106 33468 29112
rect 33692 29096 33744 29102
rect 33692 29038 33744 29044
rect 33784 29096 33836 29102
rect 33784 29038 33836 29044
rect 33704 28626 33732 29038
rect 33692 28620 33744 28626
rect 33692 28562 33744 28568
rect 33796 28490 33824 29038
rect 34348 28762 34376 29514
rect 34336 28756 34388 28762
rect 34336 28698 34388 28704
rect 33784 28484 33836 28490
rect 33784 28426 33836 28432
rect 33140 28416 33192 28422
rect 33140 28358 33192 28364
rect 33152 28150 33180 28358
rect 34334 28248 34390 28257
rect 34334 28183 34390 28192
rect 34348 28150 34376 28183
rect 34532 28150 34560 29990
rect 34624 29510 34652 30110
rect 34704 30048 34756 30054
rect 34992 30036 35020 30654
rect 35164 30592 35216 30598
rect 35164 30534 35216 30540
rect 35176 30394 35204 30534
rect 35360 30433 35388 30738
rect 35346 30424 35402 30433
rect 35164 30388 35216 30394
rect 35346 30359 35402 30368
rect 35164 30330 35216 30336
rect 35348 30320 35400 30326
rect 35348 30262 35400 30268
rect 34704 29990 34756 29996
rect 34808 30008 35020 30036
rect 34612 29504 34664 29510
rect 34612 29446 34664 29452
rect 34612 28756 34664 28762
rect 34612 28698 34664 28704
rect 33140 28144 33192 28150
rect 33140 28086 33192 28092
rect 34336 28144 34388 28150
rect 34336 28086 34388 28092
rect 34520 28144 34572 28150
rect 34520 28086 34572 28092
rect 32956 27872 33008 27878
rect 32956 27814 33008 27820
rect 32588 27668 32640 27674
rect 32588 27610 32640 27616
rect 32864 26784 32916 26790
rect 32864 26726 32916 26732
rect 32876 26586 32904 26726
rect 32312 26580 32364 26586
rect 32312 26522 32364 26528
rect 32864 26580 32916 26586
rect 32864 26522 32916 26528
rect 32968 26382 32996 27814
rect 34624 27470 34652 28698
rect 33784 27464 33836 27470
rect 33784 27406 33836 27412
rect 34612 27464 34664 27470
rect 34612 27406 34664 27412
rect 33416 27328 33468 27334
rect 33416 27270 33468 27276
rect 33428 27062 33456 27270
rect 33796 27130 33824 27406
rect 33784 27124 33836 27130
rect 33784 27066 33836 27072
rect 33416 27056 33468 27062
rect 33416 26998 33468 27004
rect 34152 27056 34204 27062
rect 34152 26998 34204 27004
rect 34164 26586 34192 26998
rect 34612 26784 34664 26790
rect 34612 26726 34664 26732
rect 34152 26580 34204 26586
rect 34152 26522 34204 26528
rect 32956 26376 33008 26382
rect 32956 26318 33008 26324
rect 31760 25288 31812 25294
rect 31760 25230 31812 25236
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 34624 24818 34652 26726
rect 34716 26450 34744 29990
rect 34808 29646 34836 30008
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35360 29850 35388 30262
rect 35452 30054 35480 33322
rect 36004 32858 36032 34904
rect 36096 33810 36124 36128
rect 36188 35494 36216 36586
rect 36176 35488 36228 35494
rect 36176 35430 36228 35436
rect 36176 35148 36228 35154
rect 36176 35090 36228 35096
rect 36188 35018 36216 35090
rect 36176 35012 36228 35018
rect 36176 34954 36228 34960
rect 36176 34400 36228 34406
rect 36176 34342 36228 34348
rect 36188 33930 36216 34342
rect 36176 33924 36228 33930
rect 36176 33866 36228 33872
rect 36096 33782 36216 33810
rect 36004 32830 36124 32858
rect 35992 32768 36044 32774
rect 35992 32710 36044 32716
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 35808 32564 35860 32570
rect 35808 32506 35860 32512
rect 35532 32428 35584 32434
rect 35532 32370 35584 32376
rect 35544 31890 35572 32370
rect 35532 31884 35584 31890
rect 35532 31826 35584 31832
rect 35820 31686 35848 32506
rect 36004 31906 36032 32710
rect 36096 32570 36124 32830
rect 36084 32564 36136 32570
rect 36084 32506 36136 32512
rect 35912 31890 36032 31906
rect 35900 31884 36032 31890
rect 35952 31878 36032 31884
rect 36084 31884 36136 31890
rect 35900 31826 35952 31832
rect 36084 31826 36136 31832
rect 35912 31754 35940 31826
rect 35912 31726 36032 31754
rect 35808 31680 35860 31686
rect 35808 31622 35860 31628
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 35808 31136 35860 31142
rect 35808 31078 35860 31084
rect 35820 30598 35848 31078
rect 35808 30592 35860 30598
rect 35808 30534 35860 30540
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 35624 30388 35676 30394
rect 35624 30330 35676 30336
rect 35440 30048 35492 30054
rect 35440 29990 35492 29996
rect 35532 30048 35584 30054
rect 35532 29990 35584 29996
rect 35348 29844 35400 29850
rect 35348 29786 35400 29792
rect 35346 29744 35402 29753
rect 35346 29679 35402 29688
rect 34796 29640 34848 29646
rect 34796 29582 34848 29588
rect 35164 29504 35216 29510
rect 35164 29446 35216 29452
rect 35256 29504 35308 29510
rect 35256 29446 35308 29452
rect 34796 29164 34848 29170
rect 34796 29106 34848 29112
rect 34808 28762 34836 29106
rect 35176 29034 35204 29446
rect 35164 29028 35216 29034
rect 35164 28970 35216 28976
rect 35268 28966 35296 29446
rect 35256 28960 35308 28966
rect 35256 28902 35308 28908
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34796 28756 34848 28762
rect 34796 28698 34848 28704
rect 34796 28552 34848 28558
rect 34796 28494 34848 28500
rect 34704 26444 34756 26450
rect 34704 26386 34756 26392
rect 34716 26042 34744 26386
rect 34808 26382 34836 28494
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35360 27062 35388 29679
rect 35544 29646 35572 29990
rect 35532 29640 35584 29646
rect 35452 29600 35532 29628
rect 35452 28558 35480 29600
rect 35532 29582 35584 29588
rect 35636 29510 35664 30330
rect 35900 30116 35952 30122
rect 35900 30058 35952 30064
rect 35912 29782 35940 30058
rect 35900 29776 35952 29782
rect 35900 29718 35952 29724
rect 36004 29578 36032 31726
rect 36096 31278 36124 31826
rect 36084 31272 36136 31278
rect 36084 31214 36136 31220
rect 36188 30666 36216 33782
rect 36280 32230 36308 43862
rect 36464 42906 36492 43948
rect 36740 43353 36768 44134
rect 37096 43988 37148 43994
rect 37096 43930 37148 43936
rect 37108 43790 37136 43930
rect 37096 43784 37148 43790
rect 37096 43726 37148 43732
rect 36726 43344 36782 43353
rect 36636 43308 36688 43314
rect 36726 43279 36728 43288
rect 36636 43250 36688 43256
rect 36780 43279 36782 43288
rect 36912 43308 36964 43314
rect 36728 43250 36780 43256
rect 36912 43250 36964 43256
rect 36452 42900 36504 42906
rect 36452 42842 36504 42848
rect 36648 42838 36676 43250
rect 36728 43104 36780 43110
rect 36728 43046 36780 43052
rect 36636 42832 36688 42838
rect 36636 42774 36688 42780
rect 36452 42356 36504 42362
rect 36452 42298 36504 42304
rect 36360 38344 36412 38350
rect 36360 38286 36412 38292
rect 36372 37874 36400 38286
rect 36360 37868 36412 37874
rect 36360 37810 36412 37816
rect 36360 37256 36412 37262
rect 36360 37198 36412 37204
rect 36372 36038 36400 37198
rect 36360 36032 36412 36038
rect 36360 35974 36412 35980
rect 36464 35578 36492 42298
rect 36648 41274 36676 42774
rect 36740 41818 36768 43046
rect 36924 42906 36952 43250
rect 37096 43104 37148 43110
rect 37096 43046 37148 43052
rect 37108 42906 37136 43046
rect 36912 42900 36964 42906
rect 36912 42842 36964 42848
rect 37096 42900 37148 42906
rect 37096 42842 37148 42848
rect 37096 42764 37148 42770
rect 37096 42706 37148 42712
rect 36728 41812 36780 41818
rect 36728 41754 36780 41760
rect 36636 41268 36688 41274
rect 36636 41210 36688 41216
rect 36636 40928 36688 40934
rect 36636 40870 36688 40876
rect 36648 40730 36676 40870
rect 36740 40730 36768 41754
rect 37108 41414 37136 42706
rect 37188 42560 37240 42566
rect 37188 42502 37240 42508
rect 37200 41546 37228 42502
rect 37188 41540 37240 41546
rect 37188 41482 37240 41488
rect 37108 41386 37228 41414
rect 36636 40724 36688 40730
rect 36636 40666 36688 40672
rect 36728 40724 36780 40730
rect 36728 40666 36780 40672
rect 37200 40594 37228 41386
rect 37292 41138 37320 44288
rect 37280 41132 37332 41138
rect 37280 41074 37332 41080
rect 37188 40588 37240 40594
rect 37188 40530 37240 40536
rect 36728 40520 36780 40526
rect 36728 40462 36780 40468
rect 37004 40520 37056 40526
rect 37004 40462 37056 40468
rect 36740 39896 36768 40462
rect 36912 39908 36964 39914
rect 36740 39868 36912 39896
rect 36544 39024 36596 39030
rect 36544 38966 36596 38972
rect 36556 38321 36584 38966
rect 36740 38486 36768 39868
rect 36912 39850 36964 39856
rect 37016 39642 37044 40462
rect 37200 40390 37228 40530
rect 37096 40384 37148 40390
rect 37096 40326 37148 40332
rect 37188 40384 37240 40390
rect 37188 40326 37240 40332
rect 37108 40050 37136 40326
rect 37096 40044 37148 40050
rect 37096 39986 37148 39992
rect 37004 39636 37056 39642
rect 37004 39578 37056 39584
rect 36912 39432 36964 39438
rect 36832 39392 36912 39420
rect 36832 38962 36860 39392
rect 36912 39374 36964 39380
rect 36912 39296 36964 39302
rect 36912 39238 36964 39244
rect 36924 38962 36952 39238
rect 36820 38956 36872 38962
rect 36820 38898 36872 38904
rect 36912 38956 36964 38962
rect 36912 38898 36964 38904
rect 36728 38480 36780 38486
rect 36728 38422 36780 38428
rect 36832 38350 36860 38898
rect 37280 38752 37332 38758
rect 37280 38694 37332 38700
rect 37292 38350 37320 38694
rect 36636 38344 36688 38350
rect 36542 38312 36598 38321
rect 36636 38286 36688 38292
rect 36820 38344 36872 38350
rect 36820 38286 36872 38292
rect 37280 38344 37332 38350
rect 37280 38286 37332 38292
rect 36542 38247 36598 38256
rect 36556 35698 36584 38247
rect 36648 37874 36676 38286
rect 36728 38208 36780 38214
rect 36728 38150 36780 38156
rect 36636 37868 36688 37874
rect 36636 37810 36688 37816
rect 36648 37398 36676 37810
rect 36636 37392 36688 37398
rect 36636 37334 36688 37340
rect 36740 37330 36768 38150
rect 36728 37324 36780 37330
rect 36728 37266 36780 37272
rect 36636 37256 36688 37262
rect 36636 37198 36688 37204
rect 36648 36922 36676 37198
rect 36636 36916 36688 36922
rect 36636 36858 36688 36864
rect 36728 36644 36780 36650
rect 36832 36632 36860 38286
rect 37188 36780 37240 36786
rect 37188 36722 37240 36728
rect 36780 36604 36860 36632
rect 36728 36586 36780 36592
rect 36636 36372 36688 36378
rect 36636 36314 36688 36320
rect 36648 36145 36676 36314
rect 36740 36242 36768 36586
rect 36728 36236 36780 36242
rect 36728 36178 36780 36184
rect 37200 36174 37228 36722
rect 37188 36168 37240 36174
rect 36634 36136 36690 36145
rect 37188 36110 37240 36116
rect 36634 36071 36690 36080
rect 37200 35894 37228 36110
rect 37200 35866 37320 35894
rect 36544 35692 36596 35698
rect 36544 35634 36596 35640
rect 36464 35550 36676 35578
rect 36360 34196 36412 34202
rect 36360 34138 36412 34144
rect 36268 32224 36320 32230
rect 36268 32166 36320 32172
rect 36280 31890 36308 32166
rect 36372 32026 36400 34138
rect 36544 34060 36596 34066
rect 36544 34002 36596 34008
rect 36556 33114 36584 34002
rect 36544 33108 36596 33114
rect 36544 33050 36596 33056
rect 36544 32360 36596 32366
rect 36544 32302 36596 32308
rect 36452 32292 36504 32298
rect 36452 32234 36504 32240
rect 36360 32020 36412 32026
rect 36360 31962 36412 31968
rect 36268 31884 36320 31890
rect 36268 31826 36320 31832
rect 36268 31680 36320 31686
rect 36268 31622 36320 31628
rect 36280 31482 36308 31622
rect 36268 31476 36320 31482
rect 36268 31418 36320 31424
rect 36464 31346 36492 32234
rect 36556 31822 36584 32302
rect 36544 31816 36596 31822
rect 36544 31758 36596 31764
rect 36452 31340 36504 31346
rect 36452 31282 36504 31288
rect 36176 30660 36228 30666
rect 36176 30602 36228 30608
rect 36360 30660 36412 30666
rect 36360 30602 36412 30608
rect 36372 30394 36400 30602
rect 36452 30592 36504 30598
rect 36452 30534 36504 30540
rect 36360 30388 36412 30394
rect 36360 30330 36412 30336
rect 36464 29850 36492 30534
rect 36452 29844 36504 29850
rect 36452 29786 36504 29792
rect 35992 29572 36044 29578
rect 35992 29514 36044 29520
rect 35624 29504 35676 29510
rect 35624 29446 35676 29452
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 36360 29232 36412 29238
rect 36358 29200 36360 29209
rect 36412 29200 36414 29209
rect 36358 29135 36414 29144
rect 36360 29096 36412 29102
rect 36360 29038 36412 29044
rect 35808 29028 35860 29034
rect 35808 28970 35860 28976
rect 35900 29028 35952 29034
rect 35900 28970 35952 28976
rect 35992 29028 36044 29034
rect 35992 28970 36044 28976
rect 35716 28960 35768 28966
rect 35716 28902 35768 28908
rect 35440 28552 35492 28558
rect 35440 28494 35492 28500
rect 35728 28422 35756 28902
rect 35820 28626 35848 28970
rect 35808 28620 35860 28626
rect 35808 28562 35860 28568
rect 35912 28558 35940 28970
rect 36004 28558 36032 28970
rect 36084 28960 36136 28966
rect 36084 28902 36136 28908
rect 35900 28552 35952 28558
rect 35900 28494 35952 28500
rect 35992 28552 36044 28558
rect 35992 28494 36044 28500
rect 36096 28490 36124 28902
rect 36372 28694 36400 29038
rect 36360 28688 36412 28694
rect 36360 28630 36412 28636
rect 36084 28484 36136 28490
rect 36084 28426 36136 28432
rect 35716 28416 35768 28422
rect 35768 28376 36032 28404
rect 35716 28358 35768 28364
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 35348 27056 35400 27062
rect 35348 26998 35400 27004
rect 36004 26994 36032 28376
rect 36648 27606 36676 35550
rect 37188 35556 37240 35562
rect 37188 35498 37240 35504
rect 37200 35154 37228 35498
rect 37188 35148 37240 35154
rect 37188 35090 37240 35096
rect 37004 35080 37056 35086
rect 37004 35022 37056 35028
rect 37016 34678 37044 35022
rect 37004 34672 37056 34678
rect 37004 34614 37056 34620
rect 37188 34536 37240 34542
rect 37188 34478 37240 34484
rect 37096 33856 37148 33862
rect 37096 33798 37148 33804
rect 37108 33454 37136 33798
rect 37096 33448 37148 33454
rect 37096 33390 37148 33396
rect 36728 33312 36780 33318
rect 36728 33254 36780 33260
rect 37096 33312 37148 33318
rect 37096 33254 37148 33260
rect 36740 33046 36768 33254
rect 36728 33040 36780 33046
rect 36728 32982 36780 32988
rect 36912 32972 36964 32978
rect 36912 32914 36964 32920
rect 36924 32366 36952 32914
rect 36912 32360 36964 32366
rect 36912 32302 36964 32308
rect 36728 31816 36780 31822
rect 36728 31758 36780 31764
rect 36740 30394 36768 31758
rect 36820 31680 36872 31686
rect 36820 31622 36872 31628
rect 36728 30388 36780 30394
rect 36728 30330 36780 30336
rect 36832 29646 36860 31622
rect 37004 31204 37056 31210
rect 37004 31146 37056 31152
rect 36820 29640 36872 29646
rect 36820 29582 36872 29588
rect 36832 29306 36860 29582
rect 36912 29572 36964 29578
rect 36912 29514 36964 29520
rect 36820 29300 36872 29306
rect 36820 29242 36872 29248
rect 36924 29170 36952 29514
rect 36912 29164 36964 29170
rect 36912 29106 36964 29112
rect 36924 28762 36952 29106
rect 36912 28756 36964 28762
rect 36912 28698 36964 28704
rect 36636 27600 36688 27606
rect 36636 27542 36688 27548
rect 36268 27532 36320 27538
rect 36268 27474 36320 27480
rect 35992 26988 36044 26994
rect 35992 26930 36044 26936
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34796 26376 34848 26382
rect 34796 26318 34848 26324
rect 35164 26308 35216 26314
rect 35164 26250 35216 26256
rect 35176 26042 35204 26250
rect 36004 26246 36032 26930
rect 36280 26926 36308 27474
rect 36636 27396 36688 27402
rect 36636 27338 36688 27344
rect 36268 26920 36320 26926
rect 36268 26862 36320 26868
rect 36176 26308 36228 26314
rect 36176 26250 36228 26256
rect 35992 26240 36044 26246
rect 35992 26182 36044 26188
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 34704 26036 34756 26042
rect 34704 25978 34756 25984
rect 35164 26036 35216 26042
rect 35164 25978 35216 25984
rect 34612 24812 34664 24818
rect 34612 24754 34664 24760
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 34716 23866 34744 25978
rect 36004 25838 36032 26182
rect 35992 25832 36044 25838
rect 35992 25774 36044 25780
rect 34796 25696 34848 25702
rect 34796 25638 34848 25644
rect 34808 25158 34836 25638
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 36188 25498 36216 26250
rect 36280 26042 36308 26862
rect 36648 26586 36676 27338
rect 36636 26580 36688 26586
rect 36636 26522 36688 26528
rect 36452 26444 36504 26450
rect 36452 26386 36504 26392
rect 36268 26036 36320 26042
rect 36268 25978 36320 25984
rect 36176 25492 36228 25498
rect 36176 25434 36228 25440
rect 36464 25294 36492 26386
rect 36544 26308 36596 26314
rect 36544 26250 36596 26256
rect 36452 25288 36504 25294
rect 36452 25230 36504 25236
rect 34796 25152 34848 25158
rect 34796 25094 34848 25100
rect 34704 23860 34756 23866
rect 34704 23802 34756 23808
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 34808 6914 34836 25094
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 36464 24954 36492 25230
rect 36556 25226 36584 26250
rect 36648 25974 36676 26522
rect 36636 25968 36688 25974
rect 36636 25910 36688 25916
rect 37016 25294 37044 31146
rect 37108 29481 37136 33254
rect 37200 32910 37228 34478
rect 37292 33522 37320 35866
rect 37384 34202 37412 46378
rect 37660 46102 37688 46514
rect 37648 46096 37700 46102
rect 37648 46038 37700 46044
rect 37556 45960 37608 45966
rect 37556 45902 37608 45908
rect 37464 45484 37516 45490
rect 37464 45426 37516 45432
rect 37476 45286 37504 45426
rect 37568 45354 37596 45902
rect 37660 45558 37688 46038
rect 37752 46034 37780 47534
rect 38108 47252 38160 47258
rect 38108 47194 38160 47200
rect 37924 47116 37976 47122
rect 37924 47058 37976 47064
rect 37832 46572 37884 46578
rect 37832 46514 37884 46520
rect 37844 46442 37872 46514
rect 37832 46436 37884 46442
rect 37832 46378 37884 46384
rect 37740 46028 37792 46034
rect 37740 45970 37792 45976
rect 37648 45552 37700 45558
rect 37648 45494 37700 45500
rect 37752 45490 37780 45970
rect 37740 45484 37792 45490
rect 37740 45426 37792 45432
rect 37832 45416 37884 45422
rect 37832 45358 37884 45364
rect 37556 45348 37608 45354
rect 37556 45290 37608 45296
rect 37464 45280 37516 45286
rect 37464 45222 37516 45228
rect 37476 44402 37504 45222
rect 37844 44878 37872 45358
rect 37832 44872 37884 44878
rect 37832 44814 37884 44820
rect 37464 44396 37516 44402
rect 37464 44338 37516 44344
rect 37476 41274 37504 44338
rect 37740 44328 37792 44334
rect 37740 44270 37792 44276
rect 37752 42548 37780 44270
rect 37844 42702 37872 44814
rect 37936 44334 37964 47058
rect 38016 46572 38068 46578
rect 38016 46514 38068 46520
rect 38028 45830 38056 46514
rect 38016 45824 38068 45830
rect 38016 45766 38068 45772
rect 38016 44940 38068 44946
rect 38016 44882 38068 44888
rect 38028 44849 38056 44882
rect 38014 44840 38070 44849
rect 38014 44775 38070 44784
rect 38120 44334 38148 47194
rect 38304 46170 38332 47942
rect 40144 47802 40172 48146
rect 40132 47796 40184 47802
rect 40132 47738 40184 47744
rect 38936 47660 38988 47666
rect 38936 47602 38988 47608
rect 38476 47184 38528 47190
rect 38476 47126 38528 47132
rect 38488 46442 38516 47126
rect 38752 46980 38804 46986
rect 38752 46922 38804 46928
rect 38568 46912 38620 46918
rect 38568 46854 38620 46860
rect 38580 46578 38608 46854
rect 38764 46714 38792 46922
rect 38948 46714 38976 47602
rect 39764 47456 39816 47462
rect 39764 47398 39816 47404
rect 39304 47048 39356 47054
rect 39304 46990 39356 46996
rect 39212 46912 39264 46918
rect 39212 46854 39264 46860
rect 38752 46708 38804 46714
rect 38752 46650 38804 46656
rect 38936 46708 38988 46714
rect 38936 46650 38988 46656
rect 38568 46572 38620 46578
rect 38568 46514 38620 46520
rect 38660 46572 38712 46578
rect 38660 46514 38712 46520
rect 38476 46436 38528 46442
rect 38476 46378 38528 46384
rect 38568 46436 38620 46442
rect 38568 46378 38620 46384
rect 38488 46170 38516 46378
rect 38292 46164 38344 46170
rect 38292 46106 38344 46112
rect 38476 46164 38528 46170
rect 38476 46106 38528 46112
rect 38304 45966 38332 46106
rect 38292 45960 38344 45966
rect 38292 45902 38344 45908
rect 38304 45082 38332 45902
rect 38292 45076 38344 45082
rect 38292 45018 38344 45024
rect 38304 44946 38332 45018
rect 38292 44940 38344 44946
rect 38292 44882 38344 44888
rect 38200 44872 38252 44878
rect 38200 44814 38252 44820
rect 38212 44402 38240 44814
rect 38200 44396 38252 44402
rect 38200 44338 38252 44344
rect 37924 44328 37976 44334
rect 37924 44270 37976 44276
rect 38108 44328 38160 44334
rect 38108 44270 38160 44276
rect 38016 44192 38068 44198
rect 38016 44134 38068 44140
rect 38028 43790 38056 44134
rect 38016 43784 38068 43790
rect 38016 43726 38068 43732
rect 38200 43716 38252 43722
rect 38200 43658 38252 43664
rect 38212 43178 38240 43658
rect 38200 43172 38252 43178
rect 38200 43114 38252 43120
rect 37924 42764 37976 42770
rect 37924 42706 37976 42712
rect 37832 42696 37884 42702
rect 37832 42638 37884 42644
rect 37752 42520 37872 42548
rect 37648 42016 37700 42022
rect 37648 41958 37700 41964
rect 37556 41676 37608 41682
rect 37556 41618 37608 41624
rect 37464 41268 37516 41274
rect 37464 41210 37516 41216
rect 37476 37466 37504 41210
rect 37568 41138 37596 41618
rect 37660 41478 37688 41958
rect 37740 41608 37792 41614
rect 37740 41550 37792 41556
rect 37648 41472 37700 41478
rect 37648 41414 37700 41420
rect 37556 41132 37608 41138
rect 37556 41074 37608 41080
rect 37568 40934 37596 41074
rect 37556 40928 37608 40934
rect 37556 40870 37608 40876
rect 37554 40760 37610 40769
rect 37554 40695 37610 40704
rect 37568 38758 37596 40695
rect 37660 40458 37688 41414
rect 37752 41002 37780 41550
rect 37740 40996 37792 41002
rect 37740 40938 37792 40944
rect 37844 40594 37872 42520
rect 37936 41614 37964 42706
rect 38016 42560 38068 42566
rect 38016 42502 38068 42508
rect 38028 42362 38056 42502
rect 38016 42356 38068 42362
rect 38016 42298 38068 42304
rect 38028 41682 38056 42298
rect 38108 42016 38160 42022
rect 38108 41958 38160 41964
rect 38016 41676 38068 41682
rect 38016 41618 38068 41624
rect 38120 41614 38148 41958
rect 37924 41608 37976 41614
rect 37924 41550 37976 41556
rect 38108 41608 38160 41614
rect 38108 41550 38160 41556
rect 37936 41414 37964 41550
rect 37936 41386 38056 41414
rect 37924 41132 37976 41138
rect 37924 41074 37976 41080
rect 37936 40730 37964 41074
rect 37924 40724 37976 40730
rect 37924 40666 37976 40672
rect 37832 40588 37884 40594
rect 37832 40530 37884 40536
rect 37648 40452 37700 40458
rect 37648 40394 37700 40400
rect 37738 40216 37794 40225
rect 37738 40151 37794 40160
rect 37752 40118 37780 40151
rect 37740 40112 37792 40118
rect 37740 40054 37792 40060
rect 37648 40044 37700 40050
rect 37648 39986 37700 39992
rect 37660 39953 37688 39986
rect 37646 39944 37702 39953
rect 37646 39879 37702 39888
rect 37660 39574 37688 39879
rect 37648 39568 37700 39574
rect 37648 39510 37700 39516
rect 37740 39568 37792 39574
rect 37740 39510 37792 39516
rect 37752 38826 37780 39510
rect 37844 39506 37872 40530
rect 37924 40452 37976 40458
rect 37924 40394 37976 40400
rect 37936 40050 37964 40394
rect 37924 40044 37976 40050
rect 37924 39986 37976 39992
rect 37832 39500 37884 39506
rect 37832 39442 37884 39448
rect 37740 38820 37792 38826
rect 37740 38762 37792 38768
rect 37556 38752 37608 38758
rect 37556 38694 37608 38700
rect 37568 37670 37596 38694
rect 37556 37664 37608 37670
rect 37556 37606 37608 37612
rect 37464 37460 37516 37466
rect 37464 37402 37516 37408
rect 37464 37120 37516 37126
rect 37464 37062 37516 37068
rect 37476 36242 37504 37062
rect 37464 36236 37516 36242
rect 37464 36178 37516 36184
rect 37476 35834 37504 36178
rect 37568 36106 37596 37606
rect 37648 37460 37700 37466
rect 37648 37402 37700 37408
rect 37660 37108 37688 37402
rect 37752 37262 37780 38762
rect 37924 38344 37976 38350
rect 37924 38286 37976 38292
rect 37832 38208 37884 38214
rect 37832 38150 37884 38156
rect 37844 37874 37872 38150
rect 37832 37868 37884 37874
rect 37832 37810 37884 37816
rect 37740 37256 37792 37262
rect 37740 37198 37792 37204
rect 37832 37120 37884 37126
rect 37660 37080 37780 37108
rect 37648 36168 37700 36174
rect 37648 36110 37700 36116
rect 37556 36100 37608 36106
rect 37556 36042 37608 36048
rect 37464 35828 37516 35834
rect 37464 35770 37516 35776
rect 37568 35698 37596 36042
rect 37464 35692 37516 35698
rect 37464 35634 37516 35640
rect 37556 35692 37608 35698
rect 37556 35634 37608 35640
rect 37476 35154 37504 35634
rect 37464 35148 37516 35154
rect 37464 35090 37516 35096
rect 37568 35034 37596 35634
rect 37660 35562 37688 36110
rect 37752 35698 37780 37080
rect 37832 37062 37884 37068
rect 37844 36854 37872 37062
rect 37832 36848 37884 36854
rect 37832 36790 37884 36796
rect 37740 35692 37792 35698
rect 37740 35634 37792 35640
rect 37648 35556 37700 35562
rect 37648 35498 37700 35504
rect 37752 35290 37780 35634
rect 37740 35284 37792 35290
rect 37740 35226 37792 35232
rect 37832 35284 37884 35290
rect 37936 35272 37964 38286
rect 38028 36718 38056 41386
rect 38108 41200 38160 41206
rect 38108 41142 38160 41148
rect 38120 40934 38148 41142
rect 38108 40928 38160 40934
rect 38108 40870 38160 40876
rect 38106 40216 38162 40225
rect 38106 40151 38108 40160
rect 38160 40151 38162 40160
rect 38108 40122 38160 40128
rect 38108 39976 38160 39982
rect 38106 39944 38108 39953
rect 38160 39944 38162 39953
rect 38106 39879 38162 39888
rect 38108 39840 38160 39846
rect 38108 39782 38160 39788
rect 38120 39506 38148 39782
rect 38108 39500 38160 39506
rect 38108 39442 38160 39448
rect 38108 38956 38160 38962
rect 38108 38898 38160 38904
rect 38120 38865 38148 38898
rect 38106 38856 38162 38865
rect 38106 38791 38162 38800
rect 38108 38344 38160 38350
rect 38106 38312 38108 38321
rect 38160 38312 38162 38321
rect 38106 38247 38162 38256
rect 38108 37460 38160 37466
rect 38108 37402 38160 37408
rect 38120 36786 38148 37402
rect 38108 36780 38160 36786
rect 38108 36722 38160 36728
rect 38016 36712 38068 36718
rect 38120 36689 38148 36722
rect 38016 36654 38068 36660
rect 38106 36680 38162 36689
rect 38106 36615 38162 36624
rect 38016 36576 38068 36582
rect 38212 36530 38240 43114
rect 38304 42022 38332 44882
rect 38384 44192 38436 44198
rect 38384 44134 38436 44140
rect 38396 43790 38424 44134
rect 38384 43784 38436 43790
rect 38384 43726 38436 43732
rect 38396 42566 38424 43726
rect 38476 43716 38528 43722
rect 38580 43704 38608 46378
rect 38672 46374 38700 46514
rect 38660 46368 38712 46374
rect 38660 46310 38712 46316
rect 38764 46102 38792 46650
rect 39224 46578 39252 46854
rect 39028 46572 39080 46578
rect 39028 46514 39080 46520
rect 39212 46572 39264 46578
rect 39212 46514 39264 46520
rect 38752 46096 38804 46102
rect 38752 46038 38804 46044
rect 38764 45948 38792 46038
rect 38844 45960 38896 45966
rect 38764 45920 38844 45948
rect 38844 45902 38896 45908
rect 38660 45892 38712 45898
rect 38660 45834 38712 45840
rect 38672 44946 38700 45834
rect 38752 45824 38804 45830
rect 38752 45766 38804 45772
rect 38660 44940 38712 44946
rect 38660 44882 38712 44888
rect 38528 43676 38608 43704
rect 38476 43658 38528 43664
rect 38384 42560 38436 42566
rect 38384 42502 38436 42508
rect 38292 42016 38344 42022
rect 38292 41958 38344 41964
rect 38384 41268 38436 41274
rect 38304 41228 38384 41256
rect 38304 39574 38332 41228
rect 38488 41256 38516 43658
rect 38672 41682 38700 44882
rect 38764 43790 38792 45766
rect 38856 44538 38884 45902
rect 39040 45830 39068 46514
rect 39028 45824 39080 45830
rect 39028 45766 39080 45772
rect 39212 45484 39264 45490
rect 39212 45426 39264 45432
rect 39224 45354 39252 45426
rect 39212 45348 39264 45354
rect 39212 45290 39264 45296
rect 38936 45280 38988 45286
rect 38936 45222 38988 45228
rect 38844 44532 38896 44538
rect 38844 44474 38896 44480
rect 38948 44402 38976 45222
rect 38936 44396 38988 44402
rect 38936 44338 38988 44344
rect 39120 44396 39172 44402
rect 39120 44338 39172 44344
rect 38752 43784 38804 43790
rect 38752 43726 38804 43732
rect 38660 41676 38712 41682
rect 38660 41618 38712 41624
rect 38436 41228 38516 41256
rect 38566 41304 38622 41313
rect 38566 41239 38568 41248
rect 38384 41210 38436 41216
rect 38620 41239 38622 41248
rect 38568 41210 38620 41216
rect 38382 41168 38438 41177
rect 38764 41138 38792 43726
rect 39132 43722 39160 44338
rect 39224 44198 39252 45290
rect 39316 45286 39344 46990
rect 39776 46578 39804 47398
rect 40040 47184 40092 47190
rect 40040 47126 40092 47132
rect 39856 47116 39908 47122
rect 39856 47058 39908 47064
rect 39764 46572 39816 46578
rect 39764 46514 39816 46520
rect 39764 45416 39816 45422
rect 39868 45404 39896 47058
rect 40052 47054 40080 47126
rect 40040 47048 40092 47054
rect 40040 46990 40092 46996
rect 39816 45376 39896 45404
rect 39764 45358 39816 45364
rect 39304 45280 39356 45286
rect 39304 45222 39356 45228
rect 39212 44192 39264 44198
rect 39212 44134 39264 44140
rect 39120 43716 39172 43722
rect 39120 43658 39172 43664
rect 38844 43648 38896 43654
rect 39028 43648 39080 43654
rect 38896 43596 39028 43602
rect 38844 43590 39080 43596
rect 38856 43574 39068 43590
rect 39316 43382 39344 45222
rect 39396 43648 39448 43654
rect 39396 43590 39448 43596
rect 39304 43376 39356 43382
rect 39210 43344 39266 43353
rect 39304 43318 39356 43324
rect 39210 43279 39212 43288
rect 39264 43279 39266 43288
rect 39212 43250 39264 43256
rect 38844 42832 38896 42838
rect 38844 42774 38896 42780
rect 38856 42158 38884 42774
rect 38936 42220 38988 42226
rect 38936 42162 38988 42168
rect 38844 42152 38896 42158
rect 38844 42094 38896 42100
rect 38948 41274 38976 42162
rect 39224 41614 39252 43250
rect 39316 43110 39344 43318
rect 39304 43104 39356 43110
rect 39304 43046 39356 43052
rect 39316 42770 39344 43046
rect 39408 42838 39436 43590
rect 39776 43246 39804 45358
rect 40144 44402 40172 47738
rect 40236 46714 40264 48690
rect 40604 48278 40632 48690
rect 40592 48272 40644 48278
rect 40592 48214 40644 48220
rect 40316 46912 40368 46918
rect 40316 46854 40368 46860
rect 40408 46912 40460 46918
rect 40408 46854 40460 46860
rect 40224 46708 40276 46714
rect 40224 46650 40276 46656
rect 40328 46578 40356 46854
rect 40316 46572 40368 46578
rect 40316 46514 40368 46520
rect 40224 46436 40276 46442
rect 40224 46378 40276 46384
rect 40236 45898 40264 46378
rect 40420 45966 40448 46854
rect 40776 46708 40828 46714
rect 40776 46650 40828 46656
rect 40684 46640 40736 46646
rect 40684 46582 40736 46588
rect 40696 46442 40724 46582
rect 40788 46442 40816 46650
rect 40684 46436 40736 46442
rect 40684 46378 40736 46384
rect 40776 46436 40828 46442
rect 40776 46378 40828 46384
rect 40500 46164 40552 46170
rect 40500 46106 40552 46112
rect 40512 45966 40540 46106
rect 40408 45960 40460 45966
rect 40408 45902 40460 45908
rect 40500 45960 40552 45966
rect 40500 45902 40552 45908
rect 40788 45948 40816 46378
rect 40868 45960 40920 45966
rect 40788 45920 40868 45948
rect 40224 45892 40276 45898
rect 40224 45834 40276 45840
rect 40236 45558 40264 45834
rect 40224 45552 40276 45558
rect 40224 45494 40276 45500
rect 40498 45520 40554 45529
rect 40132 44396 40184 44402
rect 40132 44338 40184 44344
rect 40236 43314 40264 45494
rect 40788 45490 40816 45920
rect 40868 45902 40920 45908
rect 40498 45455 40500 45464
rect 40552 45455 40554 45464
rect 40776 45484 40828 45490
rect 40500 45426 40552 45432
rect 40776 45426 40828 45432
rect 40406 43752 40462 43761
rect 40406 43687 40462 43696
rect 40420 43450 40448 43687
rect 40408 43444 40460 43450
rect 40408 43386 40460 43392
rect 40314 43344 40370 43353
rect 40040 43308 40092 43314
rect 40040 43250 40092 43256
rect 40224 43308 40276 43314
rect 40512 43330 40540 45426
rect 40684 44192 40736 44198
rect 40684 44134 40736 44140
rect 40696 43858 40724 44134
rect 40684 43852 40736 43858
rect 40684 43794 40736 43800
rect 40592 43784 40644 43790
rect 40592 43726 40644 43732
rect 40604 43450 40632 43726
rect 40592 43444 40644 43450
rect 40592 43386 40644 43392
rect 40370 43302 40540 43330
rect 40684 43308 40736 43314
rect 40314 43279 40316 43288
rect 40224 43250 40276 43256
rect 40368 43279 40370 43288
rect 40316 43250 40368 43256
rect 40788 43296 40816 45426
rect 40972 45354 41000 48690
rect 42904 48278 42932 48708
rect 43364 48618 43392 48758
rect 43352 48612 43404 48618
rect 43352 48554 43404 48560
rect 42892 48272 42944 48278
rect 42892 48214 42944 48220
rect 41236 48136 41288 48142
rect 41236 48078 41288 48084
rect 41052 46368 41104 46374
rect 41052 46310 41104 46316
rect 40960 45348 41012 45354
rect 40960 45290 41012 45296
rect 41064 45082 41092 46310
rect 41248 46170 41276 48078
rect 41788 48000 41840 48006
rect 41788 47942 41840 47948
rect 41420 47592 41472 47598
rect 41420 47534 41472 47540
rect 41328 47184 41380 47190
rect 41328 47126 41380 47132
rect 41340 46510 41368 47126
rect 41432 46714 41460 47534
rect 41512 46912 41564 46918
rect 41512 46854 41564 46860
rect 41420 46708 41472 46714
rect 41420 46650 41472 46656
rect 41328 46504 41380 46510
rect 41328 46446 41380 46452
rect 41236 46164 41288 46170
rect 41236 46106 41288 46112
rect 41052 45076 41104 45082
rect 41052 45018 41104 45024
rect 41236 44736 41288 44742
rect 41236 44678 41288 44684
rect 40868 44328 40920 44334
rect 40868 44270 40920 44276
rect 40736 43268 40816 43296
rect 40684 43250 40736 43256
rect 39488 43240 39540 43246
rect 39488 43182 39540 43188
rect 39764 43240 39816 43246
rect 39764 43182 39816 43188
rect 39396 42832 39448 42838
rect 39396 42774 39448 42780
rect 39304 42764 39356 42770
rect 39304 42706 39356 42712
rect 39304 42084 39356 42090
rect 39304 42026 39356 42032
rect 39212 41608 39264 41614
rect 39212 41550 39264 41556
rect 38936 41268 38988 41274
rect 38936 41210 38988 41216
rect 38614 41132 38666 41138
rect 38382 41103 38384 41112
rect 38436 41103 38438 41112
rect 38384 41074 38436 41080
rect 38488 41092 38614 41120
rect 38488 40730 38516 41092
rect 38614 41074 38666 41080
rect 38752 41132 38804 41138
rect 38752 41074 38804 41080
rect 38566 41032 38622 41041
rect 38566 40967 38568 40976
rect 38620 40967 38622 40976
rect 38568 40938 38620 40944
rect 38476 40724 38528 40730
rect 38476 40666 38528 40672
rect 38292 39568 38344 39574
rect 38292 39510 38344 39516
rect 38384 37324 38436 37330
rect 38488 37312 38516 40666
rect 39224 40526 39252 41550
rect 39212 40520 39264 40526
rect 39212 40462 39264 40468
rect 38568 40044 38620 40050
rect 38568 39986 38620 39992
rect 38844 40044 38896 40050
rect 38844 39986 38896 39992
rect 38436 37284 38516 37312
rect 38384 37266 38436 37272
rect 38396 36582 38424 37266
rect 38016 36518 38068 36524
rect 38028 36106 38056 36518
rect 38120 36502 38240 36530
rect 38384 36576 38436 36582
rect 38384 36518 38436 36524
rect 38016 36100 38068 36106
rect 38016 36042 38068 36048
rect 37884 35244 37964 35272
rect 37832 35226 37884 35232
rect 37476 35006 37596 35034
rect 37740 35080 37792 35086
rect 37740 35022 37792 35028
rect 37648 35012 37700 35018
rect 37372 34196 37424 34202
rect 37372 34138 37424 34144
rect 37280 33516 37332 33522
rect 37280 33458 37332 33464
rect 37188 32904 37240 32910
rect 37188 32846 37240 32852
rect 37372 32904 37424 32910
rect 37372 32846 37424 32852
rect 37200 31822 37228 32846
rect 37280 32836 37332 32842
rect 37280 32778 37332 32784
rect 37292 32609 37320 32778
rect 37278 32600 37334 32609
rect 37384 32570 37412 32846
rect 37278 32535 37334 32544
rect 37372 32564 37424 32570
rect 37372 32506 37424 32512
rect 37280 32496 37332 32502
rect 37280 32438 37332 32444
rect 37292 32026 37320 32438
rect 37280 32020 37332 32026
rect 37280 31962 37332 31968
rect 37292 31890 37320 31962
rect 37280 31884 37332 31890
rect 37280 31826 37332 31832
rect 37188 31816 37240 31822
rect 37188 31758 37240 31764
rect 37476 31226 37504 35006
rect 37648 34954 37700 34960
rect 37556 34944 37608 34950
rect 37556 34886 37608 34892
rect 37568 34066 37596 34886
rect 37660 34610 37688 34954
rect 37648 34604 37700 34610
rect 37648 34546 37700 34552
rect 37648 34400 37700 34406
rect 37648 34342 37700 34348
rect 37556 34060 37608 34066
rect 37556 34002 37608 34008
rect 37660 33930 37688 34342
rect 37648 33924 37700 33930
rect 37648 33866 37700 33872
rect 37752 33522 37780 35022
rect 37844 34542 37872 35226
rect 37832 34536 37884 34542
rect 37832 34478 37884 34484
rect 38028 33930 38056 36042
rect 37832 33924 37884 33930
rect 37832 33866 37884 33872
rect 38016 33924 38068 33930
rect 38016 33866 38068 33872
rect 37740 33516 37792 33522
rect 37740 33458 37792 33464
rect 37752 32910 37780 33458
rect 37740 32904 37792 32910
rect 37740 32846 37792 32852
rect 37648 32836 37700 32842
rect 37648 32778 37700 32784
rect 37554 32600 37610 32609
rect 37554 32535 37556 32544
rect 37608 32535 37610 32544
rect 37556 32506 37608 32512
rect 37556 32224 37608 32230
rect 37556 32166 37608 32172
rect 37568 31822 37596 32166
rect 37556 31816 37608 31822
rect 37556 31758 37608 31764
rect 37384 31198 37504 31226
rect 37280 30388 37332 30394
rect 37280 30330 37332 30336
rect 37292 29510 37320 30330
rect 37384 29714 37412 31198
rect 37464 31136 37516 31142
rect 37464 31078 37516 31084
rect 37476 30666 37504 31078
rect 37464 30660 37516 30666
rect 37464 30602 37516 30608
rect 37556 30320 37608 30326
rect 37556 30262 37608 30268
rect 37568 29782 37596 30262
rect 37556 29776 37608 29782
rect 37556 29718 37608 29724
rect 37372 29708 37424 29714
rect 37372 29650 37424 29656
rect 37280 29504 37332 29510
rect 37094 29472 37150 29481
rect 37280 29446 37332 29452
rect 37094 29407 37150 29416
rect 37292 28914 37320 29446
rect 37384 29306 37412 29650
rect 37660 29306 37688 32778
rect 37844 32065 37872 33866
rect 37924 32904 37976 32910
rect 37924 32846 37976 32852
rect 37936 32502 37964 32846
rect 37924 32496 37976 32502
rect 37924 32438 37976 32444
rect 37830 32056 37886 32065
rect 37830 31991 37886 32000
rect 38120 31482 38148 36502
rect 38292 36168 38344 36174
rect 38292 36110 38344 36116
rect 38200 35216 38252 35222
rect 38200 35158 38252 35164
rect 38212 35086 38240 35158
rect 38200 35080 38252 35086
rect 38200 35022 38252 35028
rect 38304 34610 38332 36110
rect 38384 36032 38436 36038
rect 38384 35974 38436 35980
rect 38292 34604 38344 34610
rect 38292 34546 38344 34552
rect 38200 33448 38252 33454
rect 38200 33390 38252 33396
rect 38212 32570 38240 33390
rect 38304 33318 38332 34546
rect 38292 33312 38344 33318
rect 38292 33254 38344 33260
rect 38396 32609 38424 35974
rect 38580 35698 38608 39986
rect 38856 39506 38884 39986
rect 38844 39500 38896 39506
rect 38844 39442 38896 39448
rect 38660 38956 38712 38962
rect 38660 38898 38712 38904
rect 38672 38418 38700 38898
rect 38660 38412 38712 38418
rect 38660 38354 38712 38360
rect 38936 38004 38988 38010
rect 38936 37946 38988 37952
rect 38948 36786 38976 37946
rect 39028 37324 39080 37330
rect 39028 37266 39080 37272
rect 39040 36922 39068 37266
rect 39212 37188 39264 37194
rect 39212 37130 39264 37136
rect 39224 36922 39252 37130
rect 39028 36916 39080 36922
rect 39028 36858 39080 36864
rect 39212 36916 39264 36922
rect 39212 36858 39264 36864
rect 38936 36780 38988 36786
rect 39212 36780 39264 36786
rect 38988 36740 39212 36768
rect 38936 36722 38988 36728
rect 39212 36722 39264 36728
rect 39212 36576 39264 36582
rect 39212 36518 39264 36524
rect 38660 36032 38712 36038
rect 38660 35974 38712 35980
rect 38568 35692 38620 35698
rect 38568 35634 38620 35640
rect 38672 35222 38700 35974
rect 38936 35828 38988 35834
rect 38936 35770 38988 35776
rect 38844 35760 38896 35766
rect 38844 35702 38896 35708
rect 38660 35216 38712 35222
rect 38660 35158 38712 35164
rect 38856 34950 38884 35702
rect 38948 35086 38976 35770
rect 39224 35698 39252 36518
rect 39212 35692 39264 35698
rect 39212 35634 39264 35640
rect 38936 35080 38988 35086
rect 38936 35022 38988 35028
rect 38844 34944 38896 34950
rect 38844 34886 38896 34892
rect 38660 34672 38712 34678
rect 38660 34614 38712 34620
rect 38672 34066 38700 34614
rect 38660 34060 38712 34066
rect 38660 34002 38712 34008
rect 38672 32910 38700 34002
rect 38856 33930 38884 34886
rect 39316 34785 39344 42026
rect 39302 34776 39358 34785
rect 39302 34711 39358 34720
rect 39304 34672 39356 34678
rect 39304 34614 39356 34620
rect 39120 34400 39172 34406
rect 39120 34342 39172 34348
rect 38844 33924 38896 33930
rect 38844 33866 38896 33872
rect 38856 33658 38884 33866
rect 38844 33652 38896 33658
rect 38844 33594 38896 33600
rect 38936 33584 38988 33590
rect 38936 33526 38988 33532
rect 38948 33114 38976 33526
rect 38936 33108 38988 33114
rect 38936 33050 38988 33056
rect 38568 32904 38620 32910
rect 38568 32846 38620 32852
rect 38660 32904 38712 32910
rect 38660 32846 38712 32852
rect 38580 32722 38608 32846
rect 38567 32694 38608 32722
rect 38660 32768 38712 32774
rect 38712 32728 39068 32756
rect 38660 32710 38712 32716
rect 38382 32600 38438 32609
rect 38200 32564 38252 32570
rect 38567 32586 38595 32694
rect 38567 32570 38654 32586
rect 38567 32564 38666 32570
rect 38567 32558 38614 32564
rect 38382 32535 38438 32544
rect 38200 32506 38252 32512
rect 38614 32506 38666 32512
rect 38844 32496 38896 32502
rect 38658 32464 38714 32473
rect 38476 32428 38528 32434
rect 38304 32388 38476 32416
rect 38304 31890 38332 32388
rect 38844 32438 38896 32444
rect 38658 32399 38660 32408
rect 38476 32370 38528 32376
rect 38712 32399 38714 32408
rect 38660 32370 38712 32376
rect 38382 32328 38438 32337
rect 38382 32263 38438 32272
rect 38292 31884 38344 31890
rect 38292 31826 38344 31832
rect 38108 31476 38160 31482
rect 38108 31418 38160 31424
rect 37924 30320 37976 30326
rect 37924 30262 37976 30268
rect 37832 30252 37884 30258
rect 37832 30194 37884 30200
rect 37372 29300 37424 29306
rect 37372 29242 37424 29248
rect 37648 29300 37700 29306
rect 37648 29242 37700 29248
rect 37556 29164 37608 29170
rect 37556 29106 37608 29112
rect 37292 28886 37412 28914
rect 37280 28756 37332 28762
rect 37280 28698 37332 28704
rect 37188 28620 37240 28626
rect 37188 28562 37240 28568
rect 37200 27674 37228 28562
rect 37292 27946 37320 28698
rect 37384 28422 37412 28886
rect 37568 28558 37596 29106
rect 37844 28966 37872 30194
rect 37832 28960 37884 28966
rect 37832 28902 37884 28908
rect 37556 28552 37608 28558
rect 37556 28494 37608 28500
rect 37372 28416 37424 28422
rect 37372 28358 37424 28364
rect 37384 28218 37412 28358
rect 37372 28212 37424 28218
rect 37372 28154 37424 28160
rect 37568 28082 37596 28494
rect 37936 28490 37964 30262
rect 38120 30258 38148 31418
rect 38108 30252 38160 30258
rect 38108 30194 38160 30200
rect 38200 30048 38252 30054
rect 38198 30016 38200 30025
rect 38252 30016 38254 30025
rect 38198 29951 38254 29960
rect 38108 28552 38160 28558
rect 38108 28494 38160 28500
rect 38200 28552 38252 28558
rect 38200 28494 38252 28500
rect 37924 28484 37976 28490
rect 37924 28426 37976 28432
rect 37556 28076 37608 28082
rect 37556 28018 37608 28024
rect 37280 27940 37332 27946
rect 37280 27882 37332 27888
rect 37188 27668 37240 27674
rect 37188 27610 37240 27616
rect 37200 27062 37228 27610
rect 37292 27606 37320 27882
rect 37280 27600 37332 27606
rect 37280 27542 37332 27548
rect 37188 27056 37240 27062
rect 37188 26998 37240 27004
rect 37200 26314 37228 26998
rect 37568 26858 37596 28018
rect 38120 27452 38148 28494
rect 38212 27674 38240 28494
rect 38304 28218 38332 31826
rect 38396 28626 38424 32263
rect 38658 32192 38714 32201
rect 38658 32127 38714 32136
rect 38566 32056 38622 32065
rect 38476 32020 38528 32026
rect 38672 32026 38700 32127
rect 38566 31991 38568 32000
rect 38476 31962 38528 31968
rect 38620 31991 38622 32000
rect 38660 32020 38712 32026
rect 38568 31962 38620 31968
rect 38660 31962 38712 31968
rect 38488 30054 38516 31962
rect 38856 31754 38884 32438
rect 39040 32416 39068 32728
rect 39132 32570 39160 34342
rect 39316 34202 39344 34614
rect 39304 34196 39356 34202
rect 39304 34138 39356 34144
rect 39120 32564 39172 32570
rect 39120 32506 39172 32512
rect 38948 32388 39068 32416
rect 39304 32428 39356 32434
rect 38844 31748 38896 31754
rect 38844 31690 38896 31696
rect 38856 31414 38884 31690
rect 38948 31686 38976 32388
rect 39304 32370 39356 32376
rect 39212 32360 39264 32366
rect 39212 32302 39264 32308
rect 39224 32230 39252 32302
rect 39212 32224 39264 32230
rect 39212 32166 39264 32172
rect 38936 31680 38988 31686
rect 38936 31622 38988 31628
rect 39028 31680 39080 31686
rect 39028 31622 39080 31628
rect 38844 31408 38896 31414
rect 38844 31350 38896 31356
rect 38752 31136 38804 31142
rect 38752 31078 38804 31084
rect 38764 30938 38792 31078
rect 38752 30932 38804 30938
rect 38752 30874 38804 30880
rect 38568 30320 38620 30326
rect 38568 30262 38620 30268
rect 38476 30048 38528 30054
rect 38476 29990 38528 29996
rect 38580 29782 38608 30262
rect 38660 30252 38712 30258
rect 38660 30194 38712 30200
rect 38568 29776 38620 29782
rect 38568 29718 38620 29724
rect 38672 29646 38700 30194
rect 38660 29640 38712 29646
rect 38660 29582 38712 29588
rect 38568 29096 38620 29102
rect 38568 29038 38620 29044
rect 38580 28694 38608 29038
rect 38568 28688 38620 28694
rect 38568 28630 38620 28636
rect 38384 28620 38436 28626
rect 38384 28562 38436 28568
rect 38580 28558 38608 28630
rect 38568 28552 38620 28558
rect 38568 28494 38620 28500
rect 38292 28212 38344 28218
rect 38292 28154 38344 28160
rect 38580 28014 38608 28494
rect 38672 28422 38700 29582
rect 38660 28416 38712 28422
rect 38660 28358 38712 28364
rect 38384 28008 38436 28014
rect 38384 27950 38436 27956
rect 38568 28008 38620 28014
rect 38568 27950 38620 27956
rect 38200 27668 38252 27674
rect 38200 27610 38252 27616
rect 38200 27464 38252 27470
rect 38120 27424 38200 27452
rect 38200 27406 38252 27412
rect 38212 26926 38240 27406
rect 37740 26920 37792 26926
rect 37740 26862 37792 26868
rect 38200 26920 38252 26926
rect 38200 26862 38252 26868
rect 37556 26852 37608 26858
rect 37556 26794 37608 26800
rect 37648 26376 37700 26382
rect 37752 26364 37780 26862
rect 37700 26336 37780 26364
rect 37648 26318 37700 26324
rect 37188 26308 37240 26314
rect 37188 26250 37240 26256
rect 37464 25900 37516 25906
rect 37464 25842 37516 25848
rect 37476 25498 37504 25842
rect 37464 25492 37516 25498
rect 37464 25434 37516 25440
rect 37004 25288 37056 25294
rect 37004 25230 37056 25236
rect 36544 25220 36596 25226
rect 36544 25162 36596 25168
rect 36452 24948 36504 24954
rect 36452 24890 36504 24896
rect 35992 24812 36044 24818
rect 35992 24754 36044 24760
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 36004 24410 36032 24754
rect 35992 24404 36044 24410
rect 35992 24346 36044 24352
rect 35992 24200 36044 24206
rect 35992 24142 36044 24148
rect 35072 24064 35124 24070
rect 35072 24006 35124 24012
rect 35084 23798 35112 24006
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 35072 23792 35124 23798
rect 35072 23734 35124 23740
rect 35440 23656 35492 23662
rect 35440 23598 35492 23604
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35452 23322 35480 23598
rect 35440 23316 35492 23322
rect 35440 23258 35492 23264
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35452 22098 35480 23258
rect 36004 23118 36032 24142
rect 36556 23866 36584 25162
rect 37476 24886 37504 25434
rect 37660 25362 37688 26318
rect 38016 26240 38068 26246
rect 38016 26182 38068 26188
rect 38028 25974 38056 26182
rect 38016 25968 38068 25974
rect 38016 25910 38068 25916
rect 38016 25832 38068 25838
rect 38016 25774 38068 25780
rect 38028 25498 38056 25774
rect 38108 25696 38160 25702
rect 38108 25638 38160 25644
rect 38120 25498 38148 25638
rect 38016 25492 38068 25498
rect 38016 25434 38068 25440
rect 38108 25492 38160 25498
rect 38108 25434 38160 25440
rect 37648 25356 37700 25362
rect 37648 25298 37700 25304
rect 38200 25288 38252 25294
rect 38200 25230 38252 25236
rect 37556 24948 37608 24954
rect 37556 24890 37608 24896
rect 37464 24880 37516 24886
rect 37464 24822 37516 24828
rect 37568 24614 37596 24890
rect 37832 24812 37884 24818
rect 37832 24754 37884 24760
rect 37556 24608 37608 24614
rect 37556 24550 37608 24556
rect 37372 24336 37424 24342
rect 37372 24278 37424 24284
rect 37188 24268 37240 24274
rect 37188 24210 37240 24216
rect 37200 23866 37228 24210
rect 36544 23860 36596 23866
rect 36544 23802 36596 23808
rect 37188 23860 37240 23866
rect 37188 23802 37240 23808
rect 36084 23792 36136 23798
rect 36084 23734 36136 23740
rect 36096 23254 36124 23734
rect 36084 23248 36136 23254
rect 36084 23190 36136 23196
rect 37384 23118 37412 24278
rect 35992 23112 36044 23118
rect 35992 23054 36044 23060
rect 37188 23112 37240 23118
rect 37372 23112 37424 23118
rect 37240 23060 37320 23066
rect 37188 23054 37320 23060
rect 37372 23054 37424 23060
rect 37200 23038 37320 23054
rect 37292 22982 37320 23038
rect 37280 22976 37332 22982
rect 37280 22918 37332 22924
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 37384 22642 37412 23054
rect 37568 22778 37596 24550
rect 37844 24138 37872 24754
rect 38016 24268 38068 24274
rect 38016 24210 38068 24216
rect 37832 24132 37884 24138
rect 37832 24074 37884 24080
rect 37844 23866 37872 24074
rect 37832 23860 37884 23866
rect 37832 23802 37884 23808
rect 37844 23186 37872 23802
rect 38028 23730 38056 24210
rect 38016 23724 38068 23730
rect 38016 23666 38068 23672
rect 37832 23180 37884 23186
rect 37832 23122 37884 23128
rect 37648 23044 37700 23050
rect 37648 22986 37700 22992
rect 37556 22772 37608 22778
rect 37556 22714 37608 22720
rect 37372 22636 37424 22642
rect 37372 22578 37424 22584
rect 36268 22432 36320 22438
rect 36268 22374 36320 22380
rect 36280 22234 36308 22374
rect 36268 22228 36320 22234
rect 36268 22170 36320 22176
rect 37384 22166 37412 22578
rect 37660 22438 37688 22986
rect 38028 22710 38056 23666
rect 38108 23316 38160 23322
rect 38108 23258 38160 23264
rect 38016 22704 38068 22710
rect 38016 22646 38068 22652
rect 38120 22642 38148 23258
rect 38212 22982 38240 25230
rect 38292 24676 38344 24682
rect 38292 24618 38344 24624
rect 38304 24206 38332 24618
rect 38292 24200 38344 24206
rect 38292 24142 38344 24148
rect 38396 23798 38424 27950
rect 38568 27668 38620 27674
rect 38568 27610 38620 27616
rect 38476 27328 38528 27334
rect 38476 27270 38528 27276
rect 38488 26994 38516 27270
rect 38476 26988 38528 26994
rect 38476 26930 38528 26936
rect 38580 26790 38608 27610
rect 38672 27470 38700 28358
rect 38764 27606 38792 30874
rect 38856 30598 38884 31350
rect 38948 30666 38976 31622
rect 39040 31414 39068 31622
rect 39028 31408 39080 31414
rect 39028 31350 39080 31356
rect 39040 31210 39068 31350
rect 39028 31204 39080 31210
rect 39028 31146 39080 31152
rect 38936 30660 38988 30666
rect 38936 30602 38988 30608
rect 38844 30592 38896 30598
rect 38844 30534 38896 30540
rect 38948 29714 38976 30602
rect 39040 30190 39068 31146
rect 39224 30190 39252 32166
rect 39316 31346 39344 32370
rect 39304 31340 39356 31346
rect 39304 31282 39356 31288
rect 39408 30870 39436 42774
rect 39500 41002 39528 43182
rect 39672 42764 39724 42770
rect 39672 42706 39724 42712
rect 39488 40996 39540 41002
rect 39488 40938 39540 40944
rect 39500 40458 39528 40938
rect 39684 40934 39712 42706
rect 40052 42566 40080 43250
rect 40236 42906 40264 43250
rect 40328 43219 40356 43250
rect 40316 43104 40368 43110
rect 40316 43046 40368 43052
rect 40224 42900 40276 42906
rect 40224 42842 40276 42848
rect 40040 42560 40092 42566
rect 40040 42502 40092 42508
rect 39672 40928 39724 40934
rect 39672 40870 39724 40876
rect 39488 40452 39540 40458
rect 39488 40394 39540 40400
rect 39500 38350 39528 40394
rect 39580 39432 39632 39438
rect 39580 39374 39632 39380
rect 39488 38344 39540 38350
rect 39488 38286 39540 38292
rect 39500 38010 39528 38286
rect 39592 38214 39620 39374
rect 39684 39370 39712 40870
rect 40052 40730 40080 42502
rect 40132 41608 40184 41614
rect 40224 41608 40276 41614
rect 40132 41550 40184 41556
rect 40222 41576 40224 41585
rect 40276 41576 40278 41585
rect 40144 40934 40172 41550
rect 40222 41511 40278 41520
rect 40132 40928 40184 40934
rect 40132 40870 40184 40876
rect 40040 40724 40092 40730
rect 40040 40666 40092 40672
rect 40040 40384 40092 40390
rect 40040 40326 40092 40332
rect 39856 40044 39908 40050
rect 39856 39986 39908 39992
rect 39868 39438 39896 39986
rect 39948 39568 40000 39574
rect 39946 39536 39948 39545
rect 40000 39536 40002 39545
rect 39946 39471 40002 39480
rect 39856 39432 39908 39438
rect 39856 39374 39908 39380
rect 39672 39364 39724 39370
rect 39672 39306 39724 39312
rect 39580 38208 39632 38214
rect 39580 38150 39632 38156
rect 39488 38004 39540 38010
rect 39488 37946 39540 37952
rect 39488 37868 39540 37874
rect 39488 37810 39540 37816
rect 39500 37670 39528 37810
rect 39488 37664 39540 37670
rect 39488 37606 39540 37612
rect 39500 36650 39528 37606
rect 39592 37330 39620 38150
rect 39684 37874 39712 39306
rect 39868 38894 39896 39374
rect 40052 38962 40080 40326
rect 40040 38956 40092 38962
rect 40040 38898 40092 38904
rect 39856 38888 39908 38894
rect 39856 38830 39908 38836
rect 40052 38486 40080 38898
rect 40040 38480 40092 38486
rect 40040 38422 40092 38428
rect 40132 38412 40184 38418
rect 40132 38354 40184 38360
rect 39764 38344 39816 38350
rect 39764 38286 39816 38292
rect 39776 38010 39804 38286
rect 39764 38004 39816 38010
rect 39764 37946 39816 37952
rect 39672 37868 39724 37874
rect 39672 37810 39724 37816
rect 39948 37732 40000 37738
rect 39948 37674 40000 37680
rect 39672 37392 39724 37398
rect 39672 37334 39724 37340
rect 39580 37324 39632 37330
rect 39580 37266 39632 37272
rect 39488 36644 39540 36650
rect 39488 36586 39540 36592
rect 39488 33516 39540 33522
rect 39488 33458 39540 33464
rect 39500 32910 39528 33458
rect 39488 32904 39540 32910
rect 39488 32846 39540 32852
rect 39500 31414 39528 32846
rect 39580 32428 39632 32434
rect 39580 32370 39632 32376
rect 39592 32298 39620 32370
rect 39580 32292 39632 32298
rect 39580 32234 39632 32240
rect 39488 31408 39540 31414
rect 39488 31350 39540 31356
rect 39396 30864 39448 30870
rect 39396 30806 39448 30812
rect 39028 30184 39080 30190
rect 39026 30152 39028 30161
rect 39212 30184 39264 30190
rect 39080 30152 39082 30161
rect 39212 30126 39264 30132
rect 39026 30087 39082 30096
rect 38936 29708 38988 29714
rect 38936 29650 38988 29656
rect 39040 29594 39068 30087
rect 38856 29566 39068 29594
rect 38856 29170 38884 29566
rect 38936 29504 38988 29510
rect 38936 29446 38988 29452
rect 38844 29164 38896 29170
rect 38844 29106 38896 29112
rect 38948 29102 38976 29446
rect 39210 29336 39266 29345
rect 39210 29271 39212 29280
rect 39264 29271 39266 29280
rect 39212 29242 39264 29248
rect 38936 29096 38988 29102
rect 38936 29038 38988 29044
rect 38948 28490 38976 29038
rect 39120 29028 39172 29034
rect 39224 29016 39252 29242
rect 39172 28988 39252 29016
rect 39120 28970 39172 28976
rect 38936 28484 38988 28490
rect 38936 28426 38988 28432
rect 39212 28484 39264 28490
rect 39212 28426 39264 28432
rect 38752 27600 38804 27606
rect 38752 27542 38804 27548
rect 38660 27464 38712 27470
rect 38660 27406 38712 27412
rect 38568 26784 38620 26790
rect 38568 26726 38620 26732
rect 38580 26450 38608 26726
rect 38948 26586 38976 28426
rect 39224 28082 39252 28426
rect 39500 28121 39528 31350
rect 39486 28112 39542 28121
rect 39212 28076 39264 28082
rect 39486 28047 39542 28056
rect 39212 28018 39264 28024
rect 39028 27872 39080 27878
rect 39028 27814 39080 27820
rect 39040 27538 39068 27814
rect 39028 27532 39080 27538
rect 39028 27474 39080 27480
rect 39040 27130 39068 27474
rect 39224 27402 39252 28018
rect 39488 28008 39540 28014
rect 39488 27950 39540 27956
rect 39500 27878 39528 27950
rect 39488 27872 39540 27878
rect 39488 27814 39540 27820
rect 39500 27470 39528 27814
rect 39592 27606 39620 32234
rect 39684 28694 39712 37334
rect 39960 37194 39988 37674
rect 40040 37256 40092 37262
rect 40040 37198 40092 37204
rect 39948 37188 40000 37194
rect 39948 37130 40000 37136
rect 40052 36854 40080 37198
rect 40040 36848 40092 36854
rect 40040 36790 40092 36796
rect 39948 36780 40000 36786
rect 39948 36722 40000 36728
rect 39960 36242 39988 36722
rect 39948 36236 40000 36242
rect 39948 36178 40000 36184
rect 40144 36174 40172 38354
rect 40224 38276 40276 38282
rect 40224 38218 40276 38224
rect 40236 37942 40264 38218
rect 40224 37936 40276 37942
rect 40224 37878 40276 37884
rect 40224 36780 40276 36786
rect 40224 36722 40276 36728
rect 40236 36378 40264 36722
rect 40224 36372 40276 36378
rect 40224 36314 40276 36320
rect 40132 36168 40184 36174
rect 40132 36110 40184 36116
rect 40132 36032 40184 36038
rect 40132 35974 40184 35980
rect 40144 35018 40172 35974
rect 40132 35012 40184 35018
rect 40132 34954 40184 34960
rect 40236 34066 40264 36314
rect 40328 34678 40356 43046
rect 40408 42900 40460 42906
rect 40408 42842 40460 42848
rect 40420 41546 40448 42842
rect 40696 41614 40724 43250
rect 40776 42220 40828 42226
rect 40776 42162 40828 42168
rect 40788 41818 40816 42162
rect 40776 41812 40828 41818
rect 40776 41754 40828 41760
rect 40776 41676 40828 41682
rect 40776 41618 40828 41624
rect 40684 41608 40736 41614
rect 40684 41550 40736 41556
rect 40408 41540 40460 41546
rect 40408 41482 40460 41488
rect 40420 40186 40448 41482
rect 40684 41132 40736 41138
rect 40788 41120 40816 41618
rect 40736 41092 40816 41120
rect 40684 41074 40736 41080
rect 40696 40526 40724 41074
rect 40776 40996 40828 41002
rect 40776 40938 40828 40944
rect 40788 40662 40816 40938
rect 40776 40656 40828 40662
rect 40776 40598 40828 40604
rect 40684 40520 40736 40526
rect 40684 40462 40736 40468
rect 40500 40384 40552 40390
rect 40500 40326 40552 40332
rect 40408 40180 40460 40186
rect 40408 40122 40460 40128
rect 40420 39574 40448 40122
rect 40408 39568 40460 39574
rect 40408 39510 40460 39516
rect 40408 38208 40460 38214
rect 40408 38150 40460 38156
rect 40420 37874 40448 38150
rect 40408 37868 40460 37874
rect 40408 37810 40460 37816
rect 40420 37670 40448 37810
rect 40408 37664 40460 37670
rect 40408 37606 40460 37612
rect 40512 37274 40540 40326
rect 40684 39568 40736 39574
rect 40684 39510 40736 39516
rect 40696 38350 40724 39510
rect 40684 38344 40736 38350
rect 40684 38286 40736 38292
rect 40776 38004 40828 38010
rect 40776 37946 40828 37952
rect 40788 37670 40816 37946
rect 40776 37664 40828 37670
rect 40776 37606 40828 37612
rect 40684 37392 40736 37398
rect 40684 37334 40736 37340
rect 40420 37246 40540 37274
rect 40592 37256 40644 37262
rect 40316 34672 40368 34678
rect 40316 34614 40368 34620
rect 40224 34060 40276 34066
rect 40224 34002 40276 34008
rect 39856 32972 39908 32978
rect 40420 32960 40448 37246
rect 40592 37198 40644 37204
rect 40604 36582 40632 37198
rect 40592 36576 40644 36582
rect 40592 36518 40644 36524
rect 40604 36310 40632 36518
rect 40592 36304 40644 36310
rect 40592 36246 40644 36252
rect 40696 36038 40724 37334
rect 40684 36032 40736 36038
rect 40684 35974 40736 35980
rect 39856 32914 39908 32920
rect 40144 32932 40448 32960
rect 39868 32366 39896 32914
rect 39856 32360 39908 32366
rect 39856 32302 39908 32308
rect 39868 31482 39896 32302
rect 40040 31748 40092 31754
rect 40040 31690 40092 31696
rect 39856 31476 39908 31482
rect 39856 31418 39908 31424
rect 39764 31340 39816 31346
rect 39764 31282 39816 31288
rect 39776 30734 39804 31282
rect 40052 31278 40080 31690
rect 40040 31272 40092 31278
rect 40040 31214 40092 31220
rect 39764 30728 39816 30734
rect 39764 30670 39816 30676
rect 39776 29782 39804 30670
rect 40040 30660 40092 30666
rect 40040 30602 40092 30608
rect 40052 30326 40080 30602
rect 40040 30320 40092 30326
rect 40040 30262 40092 30268
rect 39948 30252 40000 30258
rect 39948 30194 40000 30200
rect 39764 29776 39816 29782
rect 39764 29718 39816 29724
rect 39960 29170 39988 30194
rect 40052 29306 40080 30262
rect 40144 29782 40172 32932
rect 40408 32836 40460 32842
rect 40408 32778 40460 32784
rect 40420 32570 40448 32778
rect 40592 32768 40644 32774
rect 40592 32710 40644 32716
rect 40408 32564 40460 32570
rect 40408 32506 40460 32512
rect 40604 32434 40632 32710
rect 40408 32428 40460 32434
rect 40408 32370 40460 32376
rect 40592 32428 40644 32434
rect 40592 32370 40644 32376
rect 40224 32224 40276 32230
rect 40224 32166 40276 32172
rect 40236 31822 40264 32166
rect 40420 31822 40448 32370
rect 40224 31816 40276 31822
rect 40224 31758 40276 31764
rect 40408 31816 40460 31822
rect 40408 31758 40460 31764
rect 40132 29776 40184 29782
rect 40132 29718 40184 29724
rect 40132 29640 40184 29646
rect 40132 29582 40184 29588
rect 40040 29300 40092 29306
rect 40040 29242 40092 29248
rect 39948 29164 40000 29170
rect 39948 29106 40000 29112
rect 40040 28960 40092 28966
rect 40040 28902 40092 28908
rect 40052 28762 40080 28902
rect 40040 28756 40092 28762
rect 40040 28698 40092 28704
rect 39672 28688 39724 28694
rect 39672 28630 39724 28636
rect 39948 28552 40000 28558
rect 39948 28494 40000 28500
rect 39960 27674 39988 28494
rect 39948 27668 40000 27674
rect 39948 27610 40000 27616
rect 39580 27600 39632 27606
rect 39580 27542 39632 27548
rect 39488 27464 39540 27470
rect 39488 27406 39540 27412
rect 39212 27396 39264 27402
rect 39212 27338 39264 27344
rect 39028 27124 39080 27130
rect 39028 27066 39080 27072
rect 38936 26580 38988 26586
rect 38936 26522 38988 26528
rect 39224 26450 39252 27338
rect 39960 26994 39988 27610
rect 39488 26988 39540 26994
rect 39488 26930 39540 26936
rect 39948 26988 40000 26994
rect 39948 26930 40000 26936
rect 39500 26586 39528 26930
rect 39488 26580 39540 26586
rect 39488 26522 39540 26528
rect 38568 26444 38620 26450
rect 38568 26386 38620 26392
rect 39212 26444 39264 26450
rect 39212 26386 39264 26392
rect 39672 26376 39724 26382
rect 39672 26318 39724 26324
rect 39120 26036 39172 26042
rect 39120 25978 39172 25984
rect 38488 25906 38700 25922
rect 38488 25900 38712 25906
rect 38488 25894 38660 25900
rect 38488 25294 38516 25894
rect 38660 25842 38712 25848
rect 38936 25696 38988 25702
rect 38936 25638 38988 25644
rect 38476 25288 38528 25294
rect 38476 25230 38528 25236
rect 38488 24342 38516 25230
rect 38844 25220 38896 25226
rect 38844 25162 38896 25168
rect 38856 24886 38884 25162
rect 38844 24880 38896 24886
rect 38764 24828 38844 24834
rect 38764 24822 38896 24828
rect 38764 24806 38884 24822
rect 38948 24818 38976 25638
rect 39132 25498 39160 25978
rect 39120 25492 39172 25498
rect 39120 25434 39172 25440
rect 39028 25288 39080 25294
rect 39028 25230 39080 25236
rect 38936 24812 38988 24818
rect 38476 24336 38528 24342
rect 38476 24278 38528 24284
rect 38384 23792 38436 23798
rect 38384 23734 38436 23740
rect 38476 23520 38528 23526
rect 38476 23462 38528 23468
rect 38200 22976 38252 22982
rect 38200 22918 38252 22924
rect 38108 22636 38160 22642
rect 38108 22578 38160 22584
rect 38384 22568 38436 22574
rect 38384 22510 38436 22516
rect 37648 22432 37700 22438
rect 37648 22374 37700 22380
rect 37372 22160 37424 22166
rect 37372 22102 37424 22108
rect 35440 22092 35492 22098
rect 35440 22034 35492 22040
rect 37556 21956 37608 21962
rect 37556 21898 37608 21904
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 37568 21690 37596 21898
rect 37556 21684 37608 21690
rect 37556 21626 37608 21632
rect 37660 21554 37688 22374
rect 38396 21690 38424 22510
rect 38488 22030 38516 23462
rect 38568 22976 38620 22982
rect 38568 22918 38620 22924
rect 38476 22024 38528 22030
rect 38476 21966 38528 21972
rect 38580 21962 38608 22918
rect 38764 22030 38792 24806
rect 38936 24754 38988 24760
rect 38844 24744 38896 24750
rect 38844 24686 38896 24692
rect 38856 24070 38884 24686
rect 39040 24614 39068 25230
rect 39396 24812 39448 24818
rect 39396 24754 39448 24760
rect 39028 24608 39080 24614
rect 39028 24550 39080 24556
rect 39304 24608 39356 24614
rect 39304 24550 39356 24556
rect 39028 24200 39080 24206
rect 39026 24168 39028 24177
rect 39080 24168 39082 24177
rect 39026 24103 39082 24112
rect 38844 24064 38896 24070
rect 38844 24006 38896 24012
rect 38856 23118 38884 24006
rect 38844 23112 38896 23118
rect 38844 23054 38896 23060
rect 39212 23044 39264 23050
rect 39212 22986 39264 22992
rect 39120 22704 39172 22710
rect 39120 22646 39172 22652
rect 38752 22024 38804 22030
rect 38752 21966 38804 21972
rect 38568 21956 38620 21962
rect 38568 21898 38620 21904
rect 38660 21888 38712 21894
rect 38660 21830 38712 21836
rect 38384 21684 38436 21690
rect 38384 21626 38436 21632
rect 38672 21554 38700 21830
rect 39132 21690 39160 22646
rect 39224 22098 39252 22986
rect 39316 22982 39344 24550
rect 39408 23118 39436 24754
rect 39684 24682 39712 26318
rect 39856 25832 39908 25838
rect 39856 25774 39908 25780
rect 39868 25430 39896 25774
rect 39856 25424 39908 25430
rect 39856 25366 39908 25372
rect 39868 25158 39896 25366
rect 39856 25152 39908 25158
rect 39856 25094 39908 25100
rect 39672 24676 39724 24682
rect 39672 24618 39724 24624
rect 39868 24614 39896 25094
rect 39960 24750 39988 26930
rect 40052 25922 40080 28698
rect 40144 28558 40172 29582
rect 40236 28762 40264 31758
rect 40316 31476 40368 31482
rect 40316 31418 40368 31424
rect 40328 30666 40356 31418
rect 40420 30938 40448 31758
rect 40592 31408 40644 31414
rect 40592 31350 40644 31356
rect 40408 30932 40460 30938
rect 40408 30874 40460 30880
rect 40408 30728 40460 30734
rect 40408 30670 40460 30676
rect 40316 30660 40368 30666
rect 40316 30602 40368 30608
rect 40420 30546 40448 30670
rect 40500 30660 40552 30666
rect 40500 30602 40552 30608
rect 40328 30518 40448 30546
rect 40328 30122 40356 30518
rect 40512 30258 40540 30602
rect 40500 30252 40552 30258
rect 40500 30194 40552 30200
rect 40408 30184 40460 30190
rect 40408 30126 40460 30132
rect 40316 30116 40368 30122
rect 40316 30058 40368 30064
rect 40420 29889 40448 30126
rect 40406 29880 40462 29889
rect 40406 29815 40462 29824
rect 40408 29776 40460 29782
rect 40408 29718 40460 29724
rect 40316 29164 40368 29170
rect 40420 29152 40448 29718
rect 40512 29510 40540 30194
rect 40500 29504 40552 29510
rect 40500 29446 40552 29452
rect 40500 29164 40552 29170
rect 40420 29124 40500 29152
rect 40316 29106 40368 29112
rect 40500 29106 40552 29112
rect 40328 28937 40356 29106
rect 40512 29073 40540 29106
rect 40498 29064 40554 29073
rect 40498 28999 40554 29008
rect 40314 28928 40370 28937
rect 40314 28863 40370 28872
rect 40224 28756 40276 28762
rect 40224 28698 40276 28704
rect 40132 28552 40184 28558
rect 40132 28494 40184 28500
rect 40144 28014 40172 28494
rect 40328 28218 40356 28863
rect 40316 28212 40368 28218
rect 40316 28154 40368 28160
rect 40132 28008 40184 28014
rect 40132 27950 40184 27956
rect 40132 27872 40184 27878
rect 40132 27814 40184 27820
rect 40144 27674 40172 27814
rect 40132 27668 40184 27674
rect 40132 27610 40184 27616
rect 40604 27606 40632 31350
rect 40696 30326 40724 35974
rect 40788 30734 40816 37606
rect 40880 35698 40908 44270
rect 41248 44266 41276 44678
rect 41236 44260 41288 44266
rect 41236 44202 41288 44208
rect 41144 43920 41196 43926
rect 41144 43862 41196 43868
rect 40960 43648 41012 43654
rect 40960 43590 41012 43596
rect 40972 42945 41000 43590
rect 41050 43208 41106 43217
rect 41050 43143 41052 43152
rect 41104 43143 41106 43152
rect 41052 43114 41104 43120
rect 41156 43081 41184 43862
rect 41142 43072 41198 43081
rect 41142 43007 41198 43016
rect 40958 42936 41014 42945
rect 40958 42871 41014 42880
rect 40960 41608 41012 41614
rect 40960 41550 41012 41556
rect 40972 39506 41000 41550
rect 40960 39500 41012 39506
rect 40960 39442 41012 39448
rect 40972 38350 41000 39442
rect 41052 38888 41104 38894
rect 41052 38830 41104 38836
rect 41064 38554 41092 38830
rect 41052 38548 41104 38554
rect 41052 38490 41104 38496
rect 40960 38344 41012 38350
rect 40960 38286 41012 38292
rect 40868 35692 40920 35698
rect 40868 35634 40920 35640
rect 40960 35556 41012 35562
rect 40960 35498 41012 35504
rect 40868 31340 40920 31346
rect 40868 31282 40920 31288
rect 40776 30728 40828 30734
rect 40776 30670 40828 30676
rect 40880 30410 40908 31282
rect 40788 30382 40908 30410
rect 40684 30320 40736 30326
rect 40684 30262 40736 30268
rect 40684 30116 40736 30122
rect 40684 30058 40736 30064
rect 40696 28393 40724 30058
rect 40788 29238 40816 30382
rect 40868 30320 40920 30326
rect 40868 30262 40920 30268
rect 40880 30122 40908 30262
rect 40868 30116 40920 30122
rect 40868 30058 40920 30064
rect 40776 29232 40828 29238
rect 40776 29174 40828 29180
rect 40868 29232 40920 29238
rect 40972 29209 41000 35498
rect 41144 35080 41196 35086
rect 41144 35022 41196 35028
rect 41052 34740 41104 34746
rect 41052 34682 41104 34688
rect 41064 34542 41092 34682
rect 41156 34542 41184 35022
rect 41052 34536 41104 34542
rect 41052 34478 41104 34484
rect 41144 34536 41196 34542
rect 41144 34478 41196 34484
rect 41064 32978 41092 34478
rect 41052 32972 41104 32978
rect 41052 32914 41104 32920
rect 41248 32298 41276 44202
rect 41340 43994 41368 46446
rect 41524 46442 41552 46854
rect 41512 46436 41564 46442
rect 41512 46378 41564 46384
rect 41800 45898 41828 47942
rect 42524 47660 42576 47666
rect 42524 47602 42576 47608
rect 41880 47456 41932 47462
rect 41878 47424 41880 47433
rect 41932 47424 41934 47433
rect 41878 47359 41934 47368
rect 42536 47122 42564 47602
rect 42904 47598 42932 48214
rect 42892 47592 42944 47598
rect 42892 47534 42944 47540
rect 43076 47456 43128 47462
rect 43076 47398 43128 47404
rect 43088 47122 43116 47398
rect 42524 47116 42576 47122
rect 42524 47058 42576 47064
rect 43076 47116 43128 47122
rect 43076 47058 43128 47064
rect 43260 47048 43312 47054
rect 43260 46990 43312 46996
rect 42984 46912 43036 46918
rect 42984 46854 43036 46860
rect 42996 46646 43024 46854
rect 43272 46714 43300 46990
rect 43260 46708 43312 46714
rect 43260 46650 43312 46656
rect 42524 46640 42576 46646
rect 42524 46582 42576 46588
rect 42984 46640 43036 46646
rect 43364 46594 43392 48554
rect 44272 48544 44324 48550
rect 44272 48486 44324 48492
rect 44364 48544 44416 48550
rect 44364 48486 44416 48492
rect 44284 47666 44312 48486
rect 44272 47660 44324 47666
rect 44272 47602 44324 47608
rect 42984 46582 43036 46588
rect 42064 46572 42116 46578
rect 42064 46514 42116 46520
rect 41972 46436 42024 46442
rect 41972 46378 42024 46384
rect 41984 46170 42012 46378
rect 41972 46164 42024 46170
rect 41972 46106 42024 46112
rect 41788 45892 41840 45898
rect 41788 45834 41840 45840
rect 41420 45552 41472 45558
rect 41420 45494 41472 45500
rect 41432 45286 41460 45494
rect 41420 45280 41472 45286
rect 41420 45222 41472 45228
rect 41432 44538 41460 45222
rect 41420 44532 41472 44538
rect 41420 44474 41472 44480
rect 41328 43988 41380 43994
rect 41328 43930 41380 43936
rect 41340 43722 41368 43930
rect 41328 43716 41380 43722
rect 41328 43658 41380 43664
rect 41432 42378 41460 44474
rect 41512 44328 41564 44334
rect 41512 44270 41564 44276
rect 41524 43790 41552 44270
rect 41604 43852 41656 43858
rect 41604 43794 41656 43800
rect 41512 43784 41564 43790
rect 41512 43726 41564 43732
rect 41524 43330 41552 43726
rect 41616 43450 41644 43794
rect 41604 43444 41656 43450
rect 41604 43386 41656 43392
rect 41524 43302 41644 43330
rect 41800 43314 41828 45834
rect 41984 45830 42012 46106
rect 41972 45824 42024 45830
rect 41972 45766 42024 45772
rect 41984 45626 42012 45766
rect 41972 45620 42024 45626
rect 41972 45562 42024 45568
rect 41984 44878 42012 45562
rect 42076 45354 42104 46514
rect 42536 46102 42564 46582
rect 42708 46572 42760 46578
rect 42708 46514 42760 46520
rect 43076 46572 43128 46578
rect 43076 46514 43128 46520
rect 43272 46566 43392 46594
rect 43720 46640 43772 46646
rect 43720 46582 43772 46588
rect 42720 46170 42748 46514
rect 42708 46164 42760 46170
rect 43088 46152 43116 46514
rect 42708 46106 42760 46112
rect 42996 46124 43116 46152
rect 43168 46164 43220 46170
rect 42524 46096 42576 46102
rect 42524 46038 42576 46044
rect 42536 45966 42564 46038
rect 42524 45960 42576 45966
rect 42524 45902 42576 45908
rect 42800 45484 42852 45490
rect 42800 45426 42852 45432
rect 42064 45348 42116 45354
rect 42064 45290 42116 45296
rect 42812 45286 42840 45426
rect 42892 45416 42944 45422
rect 42892 45358 42944 45364
rect 42800 45280 42852 45286
rect 42800 45222 42852 45228
rect 41972 44872 42024 44878
rect 41972 44814 42024 44820
rect 42156 44872 42208 44878
rect 42156 44814 42208 44820
rect 42248 44872 42300 44878
rect 42248 44814 42300 44820
rect 42432 44872 42484 44878
rect 42432 44814 42484 44820
rect 42168 44266 42196 44814
rect 42260 44538 42288 44814
rect 42340 44804 42392 44810
rect 42340 44746 42392 44752
rect 42248 44532 42300 44538
rect 42248 44474 42300 44480
rect 42260 44402 42288 44474
rect 42248 44396 42300 44402
rect 42248 44338 42300 44344
rect 42156 44260 42208 44266
rect 42156 44202 42208 44208
rect 42156 43920 42208 43926
rect 42156 43862 42208 43868
rect 41972 43784 42024 43790
rect 41972 43726 42024 43732
rect 41512 43104 41564 43110
rect 41510 43072 41512 43081
rect 41564 43072 41566 43081
rect 41510 43007 41566 43016
rect 41616 42548 41644 43302
rect 41696 43308 41748 43314
rect 41696 43250 41748 43256
rect 41788 43308 41840 43314
rect 41788 43250 41840 43256
rect 41708 42684 41736 43250
rect 41984 43178 42012 43726
rect 42168 43217 42196 43862
rect 42352 43790 42380 44746
rect 42444 44742 42472 44814
rect 42432 44736 42484 44742
rect 42432 44678 42484 44684
rect 42432 44396 42484 44402
rect 42432 44338 42484 44344
rect 42444 44180 42472 44338
rect 42812 44180 42840 45222
rect 42904 44402 42932 45358
rect 42996 44878 43024 46124
rect 43168 46106 43220 46112
rect 43076 46028 43128 46034
rect 43076 45970 43128 45976
rect 43088 45354 43116 45970
rect 43180 45490 43208 46106
rect 43168 45484 43220 45490
rect 43168 45426 43220 45432
rect 43076 45348 43128 45354
rect 43076 45290 43128 45296
rect 43180 45082 43208 45426
rect 43168 45076 43220 45082
rect 43168 45018 43220 45024
rect 42984 44872 43036 44878
rect 42984 44814 43036 44820
rect 42892 44396 42944 44402
rect 42892 44338 42944 44344
rect 42444 44152 42840 44180
rect 42708 43988 42760 43994
rect 42708 43930 42760 43936
rect 42340 43784 42392 43790
rect 42340 43726 42392 43732
rect 42352 43450 42380 43726
rect 42524 43716 42576 43722
rect 42524 43658 42576 43664
rect 42340 43444 42392 43450
rect 42340 43386 42392 43392
rect 42536 43382 42564 43658
rect 42616 43648 42668 43654
rect 42616 43590 42668 43596
rect 42524 43376 42576 43382
rect 42524 43318 42576 43324
rect 42628 43314 42656 43590
rect 42720 43450 42748 43930
rect 42708 43444 42760 43450
rect 42708 43386 42760 43392
rect 42616 43308 42668 43314
rect 42616 43250 42668 43256
rect 42154 43208 42210 43217
rect 41972 43172 42024 43178
rect 42154 43143 42210 43152
rect 41972 43114 42024 43120
rect 41972 42900 42024 42906
rect 41972 42842 42024 42848
rect 41788 42696 41840 42702
rect 41708 42656 41788 42684
rect 41788 42638 41840 42644
rect 41696 42560 41748 42566
rect 41616 42520 41696 42548
rect 41696 42502 41748 42508
rect 41432 42350 41644 42378
rect 41512 42288 41564 42294
rect 41512 42230 41564 42236
rect 41328 41608 41380 41614
rect 41326 41576 41328 41585
rect 41380 41576 41382 41585
rect 41326 41511 41382 41520
rect 41420 39296 41472 39302
rect 41420 39238 41472 39244
rect 41432 39030 41460 39238
rect 41420 39024 41472 39030
rect 41420 38966 41472 38972
rect 41524 37262 41552 42230
rect 41512 37256 41564 37262
rect 41512 37198 41564 37204
rect 41420 36780 41472 36786
rect 41420 36722 41472 36728
rect 41432 35834 41460 36722
rect 41524 36378 41552 37198
rect 41512 36372 41564 36378
rect 41512 36314 41564 36320
rect 41512 36236 41564 36242
rect 41512 36178 41564 36184
rect 41420 35828 41472 35834
rect 41420 35770 41472 35776
rect 41524 35714 41552 36178
rect 41432 35698 41552 35714
rect 41420 35692 41552 35698
rect 41472 35686 41552 35692
rect 41420 35634 41472 35640
rect 41432 35086 41460 35634
rect 41420 35080 41472 35086
rect 41420 35022 41472 35028
rect 41512 35012 41564 35018
rect 41512 34954 41564 34960
rect 41524 33318 41552 34954
rect 41420 33312 41472 33318
rect 41420 33254 41472 33260
rect 41512 33312 41564 33318
rect 41512 33254 41564 33260
rect 41432 32842 41460 33254
rect 41420 32836 41472 32842
rect 41420 32778 41472 32784
rect 41616 32570 41644 42350
rect 41708 41138 41736 42502
rect 41800 42226 41828 42638
rect 41788 42220 41840 42226
rect 41788 42162 41840 42168
rect 41880 42220 41932 42226
rect 41880 42162 41932 42168
rect 41696 41132 41748 41138
rect 41696 41074 41748 41080
rect 41708 40526 41736 41074
rect 41696 40520 41748 40526
rect 41696 40462 41748 40468
rect 41708 40050 41736 40462
rect 41696 40044 41748 40050
rect 41696 39986 41748 39992
rect 41696 38004 41748 38010
rect 41696 37946 41748 37952
rect 41708 37738 41736 37946
rect 41696 37732 41748 37738
rect 41696 37674 41748 37680
rect 41800 37262 41828 42162
rect 41892 41682 41920 42162
rect 41880 41676 41932 41682
rect 41880 41618 41932 41624
rect 41984 41138 42012 42842
rect 42720 42702 42748 43386
rect 42812 42906 42840 44152
rect 42892 43852 42944 43858
rect 42892 43794 42944 43800
rect 42904 43382 42932 43794
rect 42996 43654 43024 44814
rect 43076 43784 43128 43790
rect 43076 43726 43128 43732
rect 42984 43648 43036 43654
rect 42984 43590 43036 43596
rect 42892 43376 42944 43382
rect 42892 43318 42944 43324
rect 42800 42900 42852 42906
rect 42800 42842 42852 42848
rect 42708 42696 42760 42702
rect 42708 42638 42760 42644
rect 42720 42294 42748 42638
rect 42708 42288 42760 42294
rect 42708 42230 42760 42236
rect 42340 42016 42392 42022
rect 42340 41958 42392 41964
rect 42352 41614 42380 41958
rect 42904 41750 42932 43318
rect 43088 43314 43116 43726
rect 43076 43308 43128 43314
rect 43076 43250 43128 43256
rect 42984 42152 43036 42158
rect 42984 42094 43036 42100
rect 42892 41744 42944 41750
rect 42892 41686 42944 41692
rect 42340 41608 42392 41614
rect 42340 41550 42392 41556
rect 42524 41608 42576 41614
rect 42524 41550 42576 41556
rect 42248 41540 42300 41546
rect 42248 41482 42300 41488
rect 41972 41132 42024 41138
rect 41972 41074 42024 41080
rect 41984 40458 42012 41074
rect 42260 40934 42288 41482
rect 42536 41206 42564 41550
rect 42340 41200 42392 41206
rect 42340 41142 42392 41148
rect 42524 41200 42576 41206
rect 42524 41142 42576 41148
rect 42352 41002 42380 41142
rect 42340 40996 42392 41002
rect 42340 40938 42392 40944
rect 42248 40928 42300 40934
rect 42248 40870 42300 40876
rect 41972 40452 42024 40458
rect 41972 40394 42024 40400
rect 41984 40118 42012 40394
rect 42064 40384 42116 40390
rect 42064 40326 42116 40332
rect 41972 40112 42024 40118
rect 41972 40054 42024 40060
rect 42076 39438 42104 40326
rect 42156 39568 42208 39574
rect 42154 39536 42156 39545
rect 42208 39536 42210 39545
rect 42154 39471 42210 39480
rect 42064 39432 42116 39438
rect 42064 39374 42116 39380
rect 41880 39364 41932 39370
rect 41880 39306 41932 39312
rect 41892 38876 41920 39306
rect 41972 38888 42024 38894
rect 41892 38848 41972 38876
rect 41892 38418 41920 38848
rect 41972 38830 42024 38836
rect 42076 38758 42104 39374
rect 42064 38752 42116 38758
rect 42064 38694 42116 38700
rect 41880 38412 41932 38418
rect 41880 38354 41932 38360
rect 41892 38010 41920 38354
rect 41880 38004 41932 38010
rect 41880 37946 41932 37952
rect 42076 37806 42104 38694
rect 42156 38208 42208 38214
rect 42156 38150 42208 38156
rect 42260 38162 42288 40870
rect 42352 40118 42380 40938
rect 42708 40656 42760 40662
rect 42708 40598 42760 40604
rect 42340 40112 42392 40118
rect 42340 40054 42392 40060
rect 42352 38282 42380 40054
rect 42524 39976 42576 39982
rect 42524 39918 42576 39924
rect 42536 39506 42564 39918
rect 42524 39500 42576 39506
rect 42524 39442 42576 39448
rect 42432 39296 42484 39302
rect 42432 39238 42484 39244
rect 42444 39030 42472 39238
rect 42432 39024 42484 39030
rect 42432 38966 42484 38972
rect 42536 38536 42564 39442
rect 42720 39438 42748 40598
rect 42708 39432 42760 39438
rect 42708 39374 42760 39380
rect 42800 39432 42852 39438
rect 42800 39374 42852 39380
rect 42812 38894 42840 39374
rect 42904 38962 42932 41686
rect 42996 41070 43024 42094
rect 43088 41546 43116 43250
rect 43076 41540 43128 41546
rect 43076 41482 43128 41488
rect 42984 41064 43036 41070
rect 42984 41006 43036 41012
rect 42996 40186 43024 41006
rect 42984 40180 43036 40186
rect 42984 40122 43036 40128
rect 42996 39370 43024 40122
rect 42984 39364 43036 39370
rect 42984 39306 43036 39312
rect 42892 38956 42944 38962
rect 42892 38898 42944 38904
rect 42800 38888 42852 38894
rect 42720 38848 42800 38876
rect 42720 38758 42748 38848
rect 42800 38830 42852 38836
rect 42708 38752 42760 38758
rect 42708 38694 42760 38700
rect 42444 38508 42564 38536
rect 42444 38282 42472 38508
rect 42524 38412 42576 38418
rect 42524 38354 42576 38360
rect 42340 38276 42392 38282
rect 42340 38218 42392 38224
rect 42432 38276 42484 38282
rect 42432 38218 42484 38224
rect 42064 37800 42116 37806
rect 42064 37742 42116 37748
rect 41972 37664 42024 37670
rect 41972 37606 42024 37612
rect 41788 37256 41840 37262
rect 41788 37198 41840 37204
rect 41800 36242 41828 37198
rect 41788 36236 41840 36242
rect 41788 36178 41840 36184
rect 41880 36168 41932 36174
rect 41880 36110 41932 36116
rect 41892 35698 41920 36110
rect 41880 35692 41932 35698
rect 41880 35634 41932 35640
rect 41892 35086 41920 35634
rect 41984 35290 42012 37606
rect 41972 35284 42024 35290
rect 41972 35226 42024 35232
rect 41880 35080 41932 35086
rect 41880 35022 41932 35028
rect 41696 34944 41748 34950
rect 41696 34886 41748 34892
rect 41708 34066 41736 34886
rect 41984 34610 42012 35226
rect 41972 34604 42024 34610
rect 41972 34546 42024 34552
rect 41696 34060 41748 34066
rect 41696 34002 41748 34008
rect 41972 33924 42024 33930
rect 41972 33866 42024 33872
rect 42064 33924 42116 33930
rect 42064 33866 42116 33872
rect 41984 33658 42012 33866
rect 41972 33652 42024 33658
rect 41972 33594 42024 33600
rect 42076 33522 42104 33866
rect 42064 33516 42116 33522
rect 42064 33458 42116 33464
rect 41878 33144 41934 33153
rect 41878 33079 41880 33088
rect 41932 33079 41934 33088
rect 41880 33050 41932 33056
rect 41604 32564 41656 32570
rect 41604 32506 41656 32512
rect 41328 32428 41380 32434
rect 41328 32370 41380 32376
rect 41236 32292 41288 32298
rect 41236 32234 41288 32240
rect 41248 32026 41276 32234
rect 41236 32020 41288 32026
rect 41236 31962 41288 31968
rect 41340 31822 41368 32370
rect 41616 32026 41644 32506
rect 41604 32020 41656 32026
rect 41604 31962 41656 31968
rect 42168 31890 42196 38150
rect 42260 38134 42472 38162
rect 42248 38004 42300 38010
rect 42248 37946 42300 37952
rect 42260 37262 42288 37946
rect 42248 37256 42300 37262
rect 42248 37198 42300 37204
rect 42340 36168 42392 36174
rect 42340 36110 42392 36116
rect 42352 35018 42380 36110
rect 42340 35012 42392 35018
rect 42340 34954 42392 34960
rect 42340 34740 42392 34746
rect 42340 34682 42392 34688
rect 42352 34066 42380 34682
rect 42340 34060 42392 34066
rect 42340 34002 42392 34008
rect 42340 32904 42392 32910
rect 42340 32846 42392 32852
rect 42156 31884 42208 31890
rect 42156 31826 42208 31832
rect 41328 31816 41380 31822
rect 41328 31758 41380 31764
rect 41340 31482 41368 31758
rect 41328 31476 41380 31482
rect 41380 31436 41460 31464
rect 41328 31418 41380 31424
rect 41328 30728 41380 30734
rect 41328 30670 41380 30676
rect 41340 30433 41368 30670
rect 41326 30424 41382 30433
rect 41052 30388 41104 30394
rect 41326 30359 41382 30368
rect 41052 30330 41104 30336
rect 41064 29753 41092 30330
rect 41328 30184 41380 30190
rect 41432 30172 41460 31436
rect 41512 31340 41564 31346
rect 41512 31282 41564 31288
rect 41524 30258 41552 31282
rect 41788 31136 41840 31142
rect 41788 31078 41840 31084
rect 41800 30666 41828 31078
rect 41788 30660 41840 30666
rect 41788 30602 41840 30608
rect 41512 30252 41564 30258
rect 41512 30194 41564 30200
rect 41380 30144 41460 30172
rect 41328 30126 41380 30132
rect 41328 29776 41380 29782
rect 41050 29744 41106 29753
rect 41328 29718 41380 29724
rect 41050 29679 41106 29688
rect 41050 29608 41106 29617
rect 41050 29543 41106 29552
rect 40868 29174 40920 29180
rect 40958 29200 41014 29209
rect 40788 29102 40816 29174
rect 40776 29096 40828 29102
rect 40776 29038 40828 29044
rect 40682 28384 40738 28393
rect 40682 28319 40738 28328
rect 40592 27600 40644 27606
rect 40592 27542 40644 27548
rect 40684 27464 40736 27470
rect 40684 27406 40736 27412
rect 40696 26994 40724 27406
rect 40788 27062 40816 29038
rect 40880 28490 40908 29174
rect 41064 29170 41092 29543
rect 41142 29336 41198 29345
rect 41142 29271 41144 29280
rect 41196 29271 41198 29280
rect 41144 29242 41196 29248
rect 40958 29135 41014 29144
rect 41052 29164 41104 29170
rect 41052 29106 41104 29112
rect 41156 28558 41184 29242
rect 41236 29164 41288 29170
rect 41236 29106 41288 29112
rect 41248 28937 41276 29106
rect 41340 28994 41368 29718
rect 41432 29238 41460 30144
rect 41524 30054 41552 30194
rect 41602 30152 41658 30161
rect 41602 30087 41658 30096
rect 41616 30054 41644 30087
rect 41512 30048 41564 30054
rect 41512 29990 41564 29996
rect 41604 30048 41656 30054
rect 41604 29990 41656 29996
rect 41510 29880 41566 29889
rect 41510 29815 41566 29824
rect 41788 29844 41840 29850
rect 41420 29232 41472 29238
rect 41420 29174 41472 29180
rect 41340 28966 41460 28994
rect 41234 28928 41290 28937
rect 41234 28863 41290 28872
rect 41432 28608 41460 28966
rect 41340 28580 41460 28608
rect 41144 28552 41196 28558
rect 41144 28494 41196 28500
rect 40868 28484 40920 28490
rect 40868 28426 40920 28432
rect 40880 27674 40908 28426
rect 41052 28416 41104 28422
rect 41052 28358 41104 28364
rect 41234 28384 41290 28393
rect 40868 27668 40920 27674
rect 40868 27610 40920 27616
rect 40776 27056 40828 27062
rect 40776 26998 40828 27004
rect 40684 26988 40736 26994
rect 40684 26930 40736 26936
rect 40224 26920 40276 26926
rect 40224 26862 40276 26868
rect 40130 26616 40186 26625
rect 40130 26551 40186 26560
rect 40144 26518 40172 26551
rect 40132 26512 40184 26518
rect 40132 26454 40184 26460
rect 40236 26450 40264 26862
rect 40224 26444 40276 26450
rect 40224 26386 40276 26392
rect 40316 26444 40368 26450
rect 40316 26386 40368 26392
rect 40052 25894 40172 25922
rect 40236 25906 40264 26386
rect 40328 26246 40356 26386
rect 40696 26382 40724 26930
rect 40500 26376 40552 26382
rect 40500 26318 40552 26324
rect 40684 26376 40736 26382
rect 40684 26318 40736 26324
rect 40316 26240 40368 26246
rect 40316 26182 40368 26188
rect 40512 25906 40540 26318
rect 40040 25764 40092 25770
rect 40040 25706 40092 25712
rect 40052 24886 40080 25706
rect 40144 25498 40172 25894
rect 40224 25900 40276 25906
rect 40224 25842 40276 25848
rect 40500 25900 40552 25906
rect 40500 25842 40552 25848
rect 40512 25498 40540 25842
rect 40132 25492 40184 25498
rect 40132 25434 40184 25440
rect 40500 25492 40552 25498
rect 40500 25434 40552 25440
rect 40144 24954 40172 25434
rect 40408 25356 40460 25362
rect 40408 25298 40460 25304
rect 40316 25152 40368 25158
rect 40316 25094 40368 25100
rect 40132 24948 40184 24954
rect 40132 24890 40184 24896
rect 40328 24886 40356 25094
rect 40040 24880 40092 24886
rect 40040 24822 40092 24828
rect 40316 24880 40368 24886
rect 40316 24822 40368 24828
rect 39948 24744 40000 24750
rect 39948 24686 40000 24692
rect 39856 24608 39908 24614
rect 39856 24550 39908 24556
rect 40052 24342 40080 24822
rect 40420 24818 40448 25298
rect 40408 24812 40460 24818
rect 40408 24754 40460 24760
rect 40040 24336 40092 24342
rect 40040 24278 40092 24284
rect 39764 24200 39816 24206
rect 39764 24142 39816 24148
rect 39856 24200 39908 24206
rect 39856 24142 39908 24148
rect 39776 23866 39804 24142
rect 39764 23860 39816 23866
rect 39764 23802 39816 23808
rect 39868 23730 39896 24142
rect 40316 24132 40368 24138
rect 40316 24074 40368 24080
rect 40328 23866 40356 24074
rect 40512 24070 40540 25434
rect 40868 25356 40920 25362
rect 40868 25298 40920 25304
rect 40880 24954 40908 25298
rect 41064 25226 41092 28358
rect 41234 28319 41290 28328
rect 41144 26988 41196 26994
rect 41144 26930 41196 26936
rect 41156 26450 41184 26930
rect 41144 26444 41196 26450
rect 41144 26386 41196 26392
rect 41156 25906 41184 26386
rect 41248 25974 41276 28319
rect 41340 27130 41368 28580
rect 41420 28484 41472 28490
rect 41420 28426 41472 28432
rect 41432 28393 41460 28426
rect 41418 28384 41474 28393
rect 41418 28319 41474 28328
rect 41420 27940 41472 27946
rect 41420 27882 41472 27888
rect 41328 27124 41380 27130
rect 41328 27066 41380 27072
rect 41340 26450 41368 27066
rect 41328 26444 41380 26450
rect 41328 26386 41380 26392
rect 41432 26042 41460 27882
rect 41524 27334 41552 29815
rect 41788 29786 41840 29792
rect 41604 29572 41656 29578
rect 41604 29514 41656 29520
rect 41696 29572 41748 29578
rect 41696 29514 41748 29520
rect 41616 28966 41644 29514
rect 41708 29306 41736 29514
rect 41696 29300 41748 29306
rect 41696 29242 41748 29248
rect 41604 28960 41656 28966
rect 41604 28902 41656 28908
rect 41616 27538 41644 28902
rect 41800 28642 41828 29786
rect 41880 29640 41932 29646
rect 41880 29582 41932 29588
rect 41892 29238 41920 29582
rect 41880 29232 41932 29238
rect 41880 29174 41932 29180
rect 41800 28614 42012 28642
rect 41788 28552 41840 28558
rect 41788 28494 41840 28500
rect 41800 28218 41828 28494
rect 41880 28484 41932 28490
rect 41880 28426 41932 28432
rect 41892 28218 41920 28426
rect 41788 28212 41840 28218
rect 41788 28154 41840 28160
rect 41880 28212 41932 28218
rect 41880 28154 41932 28160
rect 41984 28014 42012 28614
rect 42156 28416 42208 28422
rect 42156 28358 42208 28364
rect 42248 28416 42300 28422
rect 42248 28358 42300 28364
rect 41972 28008 42024 28014
rect 41972 27950 42024 27956
rect 42168 27674 42196 28358
rect 42260 28082 42288 28358
rect 42248 28076 42300 28082
rect 42248 28018 42300 28024
rect 42156 27668 42208 27674
rect 42156 27610 42208 27616
rect 41604 27532 41656 27538
rect 41604 27474 41656 27480
rect 41616 27384 41644 27474
rect 42248 27396 42300 27402
rect 41616 27356 41736 27384
rect 41512 27328 41564 27334
rect 41512 27270 41564 27276
rect 41512 26376 41564 26382
rect 41512 26318 41564 26324
rect 41420 26036 41472 26042
rect 41420 25978 41472 25984
rect 41236 25968 41288 25974
rect 41236 25910 41288 25916
rect 41144 25900 41196 25906
rect 41144 25842 41196 25848
rect 41156 25498 41184 25842
rect 41144 25492 41196 25498
rect 41144 25434 41196 25440
rect 41052 25220 41104 25226
rect 41052 25162 41104 25168
rect 40868 24948 40920 24954
rect 40868 24890 40920 24896
rect 40880 24818 40908 24890
rect 40868 24812 40920 24818
rect 40868 24754 40920 24760
rect 40960 24812 41012 24818
rect 40960 24754 41012 24760
rect 40776 24404 40828 24410
rect 40776 24346 40828 24352
rect 40500 24064 40552 24070
rect 40500 24006 40552 24012
rect 40788 23866 40816 24346
rect 40880 24206 40908 24754
rect 40972 24274 41000 24754
rect 41052 24676 41104 24682
rect 41052 24618 41104 24624
rect 40960 24268 41012 24274
rect 40960 24210 41012 24216
rect 40868 24200 40920 24206
rect 40868 24142 40920 24148
rect 41064 23866 41092 24618
rect 40316 23860 40368 23866
rect 40316 23802 40368 23808
rect 40776 23860 40828 23866
rect 40776 23802 40828 23808
rect 41052 23860 41104 23866
rect 41052 23802 41104 23808
rect 41328 23792 41380 23798
rect 41328 23734 41380 23740
rect 39856 23724 39908 23730
rect 39856 23666 39908 23672
rect 39868 23186 39896 23666
rect 41340 23526 41368 23734
rect 41328 23520 41380 23526
rect 41328 23462 41380 23468
rect 39856 23180 39908 23186
rect 39856 23122 39908 23128
rect 39396 23112 39448 23118
rect 39396 23054 39448 23060
rect 39304 22976 39356 22982
rect 39304 22918 39356 22924
rect 39868 22778 39896 23122
rect 40776 23044 40828 23050
rect 40776 22986 40828 22992
rect 40788 22778 40816 22986
rect 41524 22778 41552 26318
rect 41604 24880 41656 24886
rect 41604 24822 41656 24828
rect 41616 24614 41644 24822
rect 41708 24732 41736 27356
rect 42352 27384 42380 32846
rect 42444 31958 42472 38134
rect 42536 37806 42564 38354
rect 42800 38276 42852 38282
rect 42800 38218 42852 38224
rect 42812 38049 42840 38218
rect 42798 38040 42854 38049
rect 42798 37975 42854 37984
rect 42616 37868 42668 37874
rect 42616 37810 42668 37816
rect 42708 37868 42760 37874
rect 42708 37810 42760 37816
rect 42524 37800 42576 37806
rect 42524 37742 42576 37748
rect 42536 37126 42564 37742
rect 42628 37466 42656 37810
rect 42616 37460 42668 37466
rect 42616 37402 42668 37408
rect 42720 37194 42748 37810
rect 42708 37188 42760 37194
rect 42708 37130 42760 37136
rect 42524 37120 42576 37126
rect 42524 37062 42576 37068
rect 42524 36304 42576 36310
rect 42524 36246 42576 36252
rect 42536 34950 42564 36246
rect 42616 36168 42668 36174
rect 42616 36110 42668 36116
rect 42628 35698 42656 36110
rect 42708 36032 42760 36038
rect 42708 35974 42760 35980
rect 42720 35834 42748 35974
rect 42708 35828 42760 35834
rect 42708 35770 42760 35776
rect 42616 35692 42668 35698
rect 42616 35634 42668 35640
rect 42524 34944 42576 34950
rect 42524 34886 42576 34892
rect 42812 34524 42840 37975
rect 42904 37942 42932 38898
rect 42892 37936 42944 37942
rect 42892 37878 42944 37884
rect 42904 36786 42932 37878
rect 42892 36780 42944 36786
rect 42892 36722 42944 36728
rect 42904 36242 42932 36722
rect 42996 36718 43024 39306
rect 43088 37874 43116 41482
rect 43168 41132 43220 41138
rect 43168 41074 43220 41080
rect 43180 40050 43208 41074
rect 43168 40044 43220 40050
rect 43168 39986 43220 39992
rect 43180 39438 43208 39986
rect 43168 39432 43220 39438
rect 43168 39374 43220 39380
rect 43180 38962 43208 39374
rect 43168 38956 43220 38962
rect 43168 38898 43220 38904
rect 43076 37868 43128 37874
rect 43076 37810 43128 37816
rect 42984 36712 43036 36718
rect 42984 36654 43036 36660
rect 42984 36576 43036 36582
rect 42984 36518 43036 36524
rect 42996 36242 43024 36518
rect 42892 36236 42944 36242
rect 42892 36178 42944 36184
rect 42984 36236 43036 36242
rect 42984 36178 43036 36184
rect 43088 35834 43116 37810
rect 43272 37210 43300 46566
rect 43732 46510 43760 46582
rect 43812 46572 43864 46578
rect 43812 46514 43864 46520
rect 44180 46572 44232 46578
rect 44180 46514 44232 46520
rect 44272 46572 44324 46578
rect 44272 46514 44324 46520
rect 43720 46504 43772 46510
rect 43720 46446 43772 46452
rect 43628 45960 43680 45966
rect 43628 45902 43680 45908
rect 43640 45626 43668 45902
rect 43732 45830 43760 46446
rect 43720 45824 43772 45830
rect 43720 45766 43772 45772
rect 43628 45620 43680 45626
rect 43628 45562 43680 45568
rect 43352 44940 43404 44946
rect 43352 44882 43404 44888
rect 43364 44470 43392 44882
rect 43444 44872 43496 44878
rect 43444 44814 43496 44820
rect 43352 44464 43404 44470
rect 43352 44406 43404 44412
rect 43456 43450 43484 44814
rect 43628 44736 43680 44742
rect 43732 44724 43760 45766
rect 43824 45506 43852 46514
rect 44192 46170 44220 46514
rect 44180 46164 44232 46170
rect 44180 46106 44232 46112
rect 43996 46096 44048 46102
rect 43996 46038 44048 46044
rect 44008 45626 44036 46038
rect 44284 45966 44312 46514
rect 44272 45960 44324 45966
rect 44272 45902 44324 45908
rect 43996 45620 44048 45626
rect 43996 45562 44048 45568
rect 43824 45478 43944 45506
rect 43812 45416 43864 45422
rect 43812 45358 43864 45364
rect 43824 45082 43852 45358
rect 43916 45354 43944 45478
rect 43904 45348 43956 45354
rect 43904 45290 43956 45296
rect 43812 45076 43864 45082
rect 43812 45018 43864 45024
rect 44008 44962 44036 45562
rect 43680 44696 43760 44724
rect 43916 44934 44036 44962
rect 43628 44678 43680 44684
rect 43536 44328 43588 44334
rect 43536 44270 43588 44276
rect 43548 43994 43576 44270
rect 43536 43988 43588 43994
rect 43536 43930 43588 43936
rect 43444 43444 43496 43450
rect 43444 43386 43496 43392
rect 43640 43382 43668 44678
rect 43916 44538 43944 44934
rect 43996 44872 44048 44878
rect 43996 44814 44048 44820
rect 43904 44532 43956 44538
rect 43904 44474 43956 44480
rect 44008 44334 44036 44814
rect 43996 44328 44048 44334
rect 43996 44270 44048 44276
rect 43812 43988 43864 43994
rect 43812 43930 43864 43936
rect 43628 43376 43680 43382
rect 43628 43318 43680 43324
rect 43444 42900 43496 42906
rect 43444 42842 43496 42848
rect 43456 42702 43484 42842
rect 43444 42696 43496 42702
rect 43444 42638 43496 42644
rect 43352 42560 43404 42566
rect 43352 42502 43404 42508
rect 43364 42226 43392 42502
rect 43640 42226 43668 43318
rect 43720 43308 43772 43314
rect 43720 43250 43772 43256
rect 43732 43178 43760 43250
rect 43720 43172 43772 43178
rect 43720 43114 43772 43120
rect 43824 42838 43852 43930
rect 44272 43716 44324 43722
rect 44272 43658 44324 43664
rect 44180 43648 44232 43654
rect 44180 43590 44232 43596
rect 44192 43314 44220 43590
rect 44284 43382 44312 43658
rect 44272 43376 44324 43382
rect 44272 43318 44324 43324
rect 43904 43308 43956 43314
rect 44180 43308 44232 43314
rect 43904 43250 43956 43256
rect 44008 43268 44180 43296
rect 43812 42832 43864 42838
rect 43812 42774 43864 42780
rect 43916 42702 43944 43250
rect 43904 42696 43956 42702
rect 43904 42638 43956 42644
rect 43720 42560 43772 42566
rect 43720 42502 43772 42508
rect 43352 42220 43404 42226
rect 43352 42162 43404 42168
rect 43536 42220 43588 42226
rect 43536 42162 43588 42168
rect 43628 42220 43680 42226
rect 43628 42162 43680 42168
rect 43548 42106 43576 42162
rect 43732 42106 43760 42502
rect 43904 42220 43956 42226
rect 44008 42208 44036 43268
rect 44180 43250 44232 43256
rect 44180 43172 44232 43178
rect 44180 43114 44232 43120
rect 44192 42634 44220 43114
rect 44284 42770 44312 43318
rect 44376 43246 44404 48486
rect 44456 47660 44508 47666
rect 44456 47602 44508 47608
rect 46480 47660 46532 47666
rect 46480 47602 46532 47608
rect 44468 46170 44496 47602
rect 45836 47592 45888 47598
rect 45836 47534 45888 47540
rect 46388 47592 46440 47598
rect 46388 47534 46440 47540
rect 45008 47184 45060 47190
rect 45008 47126 45060 47132
rect 44640 46912 44692 46918
rect 44640 46854 44692 46860
rect 44652 46442 44680 46854
rect 45020 46578 45048 47126
rect 45848 47122 45876 47534
rect 46400 47190 46428 47534
rect 46388 47184 46440 47190
rect 46388 47126 46440 47132
rect 45836 47116 45888 47122
rect 45836 47058 45888 47064
rect 45376 47048 45428 47054
rect 45376 46990 45428 46996
rect 45388 46714 45416 46990
rect 45376 46708 45428 46714
rect 45376 46650 45428 46656
rect 45008 46572 45060 46578
rect 45008 46514 45060 46520
rect 45100 46572 45152 46578
rect 45100 46514 45152 46520
rect 45112 46458 45140 46514
rect 44640 46436 44692 46442
rect 44640 46378 44692 46384
rect 45020 46430 45140 46458
rect 44456 46164 44508 46170
rect 44456 46106 44508 46112
rect 44640 45892 44692 45898
rect 44640 45834 44692 45840
rect 44652 45529 44680 45834
rect 44638 45520 44694 45529
rect 45020 45490 45048 46430
rect 44638 45455 44694 45464
rect 45008 45484 45060 45490
rect 44456 44736 44508 44742
rect 44456 44678 44508 44684
rect 44468 44470 44496 44678
rect 44456 44464 44508 44470
rect 44456 44406 44508 44412
rect 44364 43240 44416 43246
rect 44364 43182 44416 43188
rect 44272 42764 44324 42770
rect 44272 42706 44324 42712
rect 44364 42696 44416 42702
rect 44364 42638 44416 42644
rect 44180 42628 44232 42634
rect 44180 42570 44232 42576
rect 44272 42628 44324 42634
rect 44272 42570 44324 42576
rect 44284 42362 44312 42570
rect 44272 42356 44324 42362
rect 44272 42298 44324 42304
rect 43956 42180 44036 42208
rect 43904 42162 43956 42168
rect 43548 42078 43760 42106
rect 43732 41478 43760 42078
rect 43904 41676 43956 41682
rect 43904 41618 43956 41624
rect 43720 41472 43772 41478
rect 43720 41414 43772 41420
rect 43916 41138 43944 41618
rect 44008 41206 44036 42180
rect 44272 42016 44324 42022
rect 44376 42004 44404 42638
rect 44324 41976 44404 42004
rect 44272 41958 44324 41964
rect 44284 41274 44312 41958
rect 44272 41268 44324 41274
rect 44272 41210 44324 41216
rect 43996 41200 44048 41206
rect 43996 41142 44048 41148
rect 43904 41132 43956 41138
rect 43904 41074 43956 41080
rect 43536 39976 43588 39982
rect 43536 39918 43588 39924
rect 43548 38350 43576 39918
rect 43916 39846 43944 41074
rect 44468 40050 44496 44406
rect 44548 43648 44600 43654
rect 44548 43590 44600 43596
rect 44560 42702 44588 43590
rect 44652 42838 44680 45455
rect 45008 45426 45060 45432
rect 45100 45484 45152 45490
rect 45100 45426 45152 45432
rect 45020 44810 45048 45426
rect 45112 45014 45140 45426
rect 45744 45416 45796 45422
rect 45744 45358 45796 45364
rect 45100 45008 45152 45014
rect 45100 44950 45152 44956
rect 45376 44872 45428 44878
rect 45376 44814 45428 44820
rect 45008 44804 45060 44810
rect 45008 44746 45060 44752
rect 45284 43852 45336 43858
rect 45284 43794 45336 43800
rect 44640 42832 44692 42838
rect 44640 42774 44692 42780
rect 45008 42764 45060 42770
rect 45008 42706 45060 42712
rect 44548 42696 44600 42702
rect 44548 42638 44600 42644
rect 45020 41290 45048 42706
rect 45296 42226 45324 43794
rect 45388 43790 45416 44814
rect 45756 43926 45784 45358
rect 45744 43920 45796 43926
rect 45744 43862 45796 43868
rect 45376 43784 45428 43790
rect 45374 43752 45376 43761
rect 45428 43752 45430 43761
rect 45374 43687 45430 43696
rect 45376 43172 45428 43178
rect 45376 43114 45428 43120
rect 45284 42220 45336 42226
rect 45284 42162 45336 42168
rect 45100 42152 45152 42158
rect 45100 42094 45152 42100
rect 45112 41818 45140 42094
rect 45100 41812 45152 41818
rect 45100 41754 45152 41760
rect 45020 41262 45140 41290
rect 45008 40724 45060 40730
rect 45112 40712 45140 41262
rect 45060 40684 45140 40712
rect 45008 40666 45060 40672
rect 44456 40044 44508 40050
rect 44456 39986 44508 39992
rect 43904 39840 43956 39846
rect 43904 39782 43956 39788
rect 44272 39432 44324 39438
rect 44272 39374 44324 39380
rect 44284 39098 44312 39374
rect 44272 39092 44324 39098
rect 44272 39034 44324 39040
rect 44180 38956 44232 38962
rect 44180 38898 44232 38904
rect 45008 38956 45060 38962
rect 45008 38898 45060 38904
rect 43812 38752 43864 38758
rect 43812 38694 43864 38700
rect 43536 38344 43588 38350
rect 43536 38286 43588 38292
rect 43352 37664 43404 37670
rect 43352 37606 43404 37612
rect 43364 37330 43392 37606
rect 43352 37324 43404 37330
rect 43352 37266 43404 37272
rect 43444 37256 43496 37262
rect 43272 37182 43392 37210
rect 43444 37198 43496 37204
rect 43168 36168 43220 36174
rect 43168 36110 43220 36116
rect 43076 35828 43128 35834
rect 43076 35770 43128 35776
rect 43180 35698 43208 36110
rect 43168 35692 43220 35698
rect 43168 35634 43220 35640
rect 43180 35086 43208 35634
rect 43260 35148 43312 35154
rect 43260 35090 43312 35096
rect 43168 35080 43220 35086
rect 43168 35022 43220 35028
rect 42984 35012 43036 35018
rect 42984 34954 43036 34960
rect 42536 34496 42840 34524
rect 42432 31952 42484 31958
rect 42432 31894 42484 31900
rect 42444 31210 42472 31894
rect 42432 31204 42484 31210
rect 42432 31146 42484 31152
rect 42536 29510 42564 34496
rect 42996 34066 43024 34954
rect 43168 34604 43220 34610
rect 43168 34546 43220 34552
rect 43180 34082 43208 34546
rect 43272 34202 43300 35090
rect 43260 34196 43312 34202
rect 43260 34138 43312 34144
rect 42984 34060 43036 34066
rect 43180 34054 43300 34082
rect 42984 34002 43036 34008
rect 43168 33992 43220 33998
rect 43168 33934 43220 33940
rect 42616 33924 42668 33930
rect 42616 33866 42668 33872
rect 42524 29504 42576 29510
rect 42524 29446 42576 29452
rect 42522 28112 42578 28121
rect 42522 28047 42524 28056
rect 42576 28047 42578 28056
rect 42524 28018 42576 28024
rect 42300 27356 42380 27384
rect 42248 27338 42300 27344
rect 42536 27062 42564 28018
rect 42524 27056 42576 27062
rect 42524 26998 42576 27004
rect 42432 26920 42484 26926
rect 42432 26862 42484 26868
rect 42444 26518 42472 26862
rect 42432 26512 42484 26518
rect 42432 26454 42484 26460
rect 42628 26042 42656 33866
rect 42800 33856 42852 33862
rect 42800 33798 42852 33804
rect 42708 33448 42760 33454
rect 42708 33390 42760 33396
rect 42720 32910 42748 33390
rect 42708 32904 42760 32910
rect 42708 32846 42760 32852
rect 42812 32858 42840 33798
rect 43180 33454 43208 33934
rect 43272 33862 43300 34054
rect 43364 33998 43392 37182
rect 43456 34354 43484 37198
rect 43548 36922 43576 38286
rect 43824 37942 43852 38694
rect 44192 38486 44220 38898
rect 44180 38480 44232 38486
rect 44180 38422 44232 38428
rect 43812 37936 43864 37942
rect 43812 37878 43864 37884
rect 43720 37800 43772 37806
rect 43720 37742 43772 37748
rect 43732 37466 43760 37742
rect 43720 37460 43772 37466
rect 43720 37402 43772 37408
rect 45020 37126 45048 38898
rect 45112 37126 45140 40684
rect 45284 40588 45336 40594
rect 45284 40530 45336 40536
rect 45192 40452 45244 40458
rect 45192 40394 45244 40400
rect 45204 38962 45232 40394
rect 45296 40186 45324 40530
rect 45284 40180 45336 40186
rect 45284 40122 45336 40128
rect 45192 38956 45244 38962
rect 45192 38898 45244 38904
rect 45284 37936 45336 37942
rect 45284 37878 45336 37884
rect 45008 37120 45060 37126
rect 45008 37062 45060 37068
rect 45100 37120 45152 37126
rect 45100 37062 45152 37068
rect 43536 36916 43588 36922
rect 43536 36858 43588 36864
rect 44088 36848 44140 36854
rect 44088 36790 44140 36796
rect 43996 36576 44048 36582
rect 43996 36518 44048 36524
rect 43536 35216 43588 35222
rect 43536 35158 43588 35164
rect 43548 34542 43576 35158
rect 44008 35086 44036 36518
rect 44100 35698 44128 36790
rect 44272 36780 44324 36786
rect 44272 36722 44324 36728
rect 44180 36712 44232 36718
rect 44180 36654 44232 36660
rect 44192 35698 44220 36654
rect 44284 36038 44312 36722
rect 44916 36304 44968 36310
rect 44916 36246 44968 36252
rect 44456 36168 44508 36174
rect 44456 36110 44508 36116
rect 44272 36032 44324 36038
rect 44272 35974 44324 35980
rect 44088 35692 44140 35698
rect 44088 35634 44140 35640
rect 44180 35692 44232 35698
rect 44180 35634 44232 35640
rect 44100 35562 44128 35634
rect 44088 35556 44140 35562
rect 44088 35498 44140 35504
rect 43996 35080 44048 35086
rect 43996 35022 44048 35028
rect 43904 34944 43956 34950
rect 43904 34886 43956 34892
rect 43810 34776 43866 34785
rect 43720 34740 43772 34746
rect 43810 34711 43866 34720
rect 43720 34682 43772 34688
rect 43536 34536 43588 34542
rect 43536 34478 43588 34484
rect 43456 34326 43576 34354
rect 43352 33992 43404 33998
rect 43352 33934 43404 33940
rect 43260 33856 43312 33862
rect 43260 33798 43312 33804
rect 43168 33448 43220 33454
rect 43168 33390 43220 33396
rect 42984 33380 43036 33386
rect 42984 33322 43036 33328
rect 42812 32830 42932 32858
rect 42800 32768 42852 32774
rect 42800 32710 42852 32716
rect 42812 32434 42840 32710
rect 42904 32570 42932 32830
rect 42892 32564 42944 32570
rect 42892 32506 42944 32512
rect 42800 32428 42852 32434
rect 42800 32370 42852 32376
rect 42812 31822 42840 32370
rect 42904 32026 42932 32506
rect 42996 32434 43024 33322
rect 43076 32836 43128 32842
rect 43180 32824 43208 33390
rect 43128 32796 43208 32824
rect 43076 32778 43128 32784
rect 42984 32428 43036 32434
rect 43036 32388 43116 32416
rect 42984 32370 43036 32376
rect 42892 32020 42944 32026
rect 42892 31962 42944 31968
rect 42892 31884 42944 31890
rect 42892 31826 42944 31832
rect 42800 31816 42852 31822
rect 42800 31758 42852 31764
rect 42904 31754 42932 31826
rect 43088 31822 43116 32388
rect 43076 31816 43128 31822
rect 43076 31758 43128 31764
rect 43180 31770 43208 32796
rect 43272 31890 43300 33798
rect 43352 33516 43404 33522
rect 43352 33458 43404 33464
rect 43364 32910 43392 33458
rect 43352 32904 43404 32910
rect 43352 32846 43404 32852
rect 43548 32842 43576 34326
rect 43628 34060 43680 34066
rect 43628 34002 43680 34008
rect 43536 32836 43588 32842
rect 43536 32778 43588 32784
rect 43260 31884 43312 31890
rect 43260 31826 43312 31832
rect 42892 31748 42944 31754
rect 43180 31742 43300 31770
rect 42892 31690 42944 31696
rect 42904 31278 42932 31690
rect 43076 31680 43128 31686
rect 43076 31622 43128 31628
rect 42892 31272 42944 31278
rect 42706 31240 42762 31249
rect 42892 31214 42944 31220
rect 42984 31272 43036 31278
rect 42984 31214 43036 31220
rect 42706 31175 42708 31184
rect 42760 31175 42762 31184
rect 42708 31146 42760 31152
rect 42720 29850 42748 31146
rect 42800 30252 42852 30258
rect 42800 30194 42852 30200
rect 42708 29844 42760 29850
rect 42708 29786 42760 29792
rect 42706 29744 42762 29753
rect 42812 29714 42840 30194
rect 42996 30122 43024 31214
rect 43088 30734 43116 31622
rect 43168 31204 43220 31210
rect 43168 31146 43220 31152
rect 43076 30728 43128 30734
rect 43076 30670 43128 30676
rect 43180 30258 43208 31146
rect 43168 30252 43220 30258
rect 43168 30194 43220 30200
rect 42984 30116 43036 30122
rect 42984 30058 43036 30064
rect 42982 30016 43038 30025
rect 42982 29951 43038 29960
rect 42706 29679 42762 29688
rect 42800 29708 42852 29714
rect 42720 28966 42748 29679
rect 42800 29650 42852 29656
rect 42708 28960 42760 28966
rect 42708 28902 42760 28908
rect 42720 28626 42748 28902
rect 42708 28620 42760 28626
rect 42708 28562 42760 28568
rect 42812 27554 42840 29650
rect 42996 29170 43024 29951
rect 43076 29504 43128 29510
rect 43076 29446 43128 29452
rect 42984 29164 43036 29170
rect 42984 29106 43036 29112
rect 42984 27872 43036 27878
rect 42984 27814 43036 27820
rect 42720 27538 42840 27554
rect 42708 27532 42840 27538
rect 42760 27526 42840 27532
rect 42708 27474 42760 27480
rect 42720 26450 42748 27474
rect 42996 27402 43024 27814
rect 42984 27396 43036 27402
rect 42984 27338 43036 27344
rect 42984 26988 43036 26994
rect 42984 26930 43036 26936
rect 42708 26444 42760 26450
rect 42708 26386 42760 26392
rect 42248 26036 42300 26042
rect 42248 25978 42300 25984
rect 42616 26036 42668 26042
rect 42616 25978 42668 25984
rect 41972 25900 42024 25906
rect 41972 25842 42024 25848
rect 41984 24818 42012 25842
rect 42260 25158 42288 25978
rect 42720 25362 42748 26386
rect 42996 25906 43024 26930
rect 42984 25900 43036 25906
rect 42984 25842 43036 25848
rect 42708 25356 42760 25362
rect 42708 25298 42760 25304
rect 42248 25152 42300 25158
rect 42248 25094 42300 25100
rect 41972 24812 42024 24818
rect 41972 24754 42024 24760
rect 42720 24750 42748 25298
rect 42892 24812 42944 24818
rect 42892 24754 42944 24760
rect 41788 24744 41840 24750
rect 41708 24704 41788 24732
rect 41788 24686 41840 24692
rect 42708 24744 42760 24750
rect 42708 24686 42760 24692
rect 41604 24608 41656 24614
rect 41604 24550 41656 24556
rect 41604 24200 41656 24206
rect 41602 24168 41604 24177
rect 41656 24168 41658 24177
rect 41602 24103 41658 24112
rect 41800 23322 41828 24686
rect 42156 24132 42208 24138
rect 42156 24074 42208 24080
rect 42064 23724 42116 23730
rect 42064 23666 42116 23672
rect 41788 23316 41840 23322
rect 41788 23258 41840 23264
rect 42076 23186 42104 23666
rect 42064 23180 42116 23186
rect 42064 23122 42116 23128
rect 42168 23050 42196 24074
rect 42720 23730 42748 24686
rect 42904 24206 42932 24754
rect 42892 24200 42944 24206
rect 42892 24142 42944 24148
rect 42708 23724 42760 23730
rect 42708 23666 42760 23672
rect 42156 23044 42208 23050
rect 42156 22986 42208 22992
rect 39856 22772 39908 22778
rect 39856 22714 39908 22720
rect 40776 22772 40828 22778
rect 40776 22714 40828 22720
rect 41512 22772 41564 22778
rect 41512 22714 41564 22720
rect 42720 22642 42748 23666
rect 42996 23526 43024 25842
rect 43088 25498 43116 29446
rect 43272 28558 43300 31742
rect 43352 31340 43404 31346
rect 43352 31282 43404 31288
rect 43364 30802 43392 31282
rect 43444 31136 43496 31142
rect 43444 31078 43496 31084
rect 43352 30796 43404 30802
rect 43352 30738 43404 30744
rect 43456 30666 43484 31078
rect 43444 30660 43496 30666
rect 43444 30602 43496 30608
rect 43352 29640 43404 29646
rect 43352 29582 43404 29588
rect 43364 29306 43392 29582
rect 43352 29300 43404 29306
rect 43352 29242 43404 29248
rect 43260 28552 43312 28558
rect 43260 28494 43312 28500
rect 43168 28212 43220 28218
rect 43168 28154 43220 28160
rect 43076 25492 43128 25498
rect 43076 25434 43128 25440
rect 43180 25430 43208 28154
rect 43272 27674 43300 28494
rect 43260 27668 43312 27674
rect 43260 27610 43312 27616
rect 43640 26790 43668 34002
rect 43732 32570 43760 34682
rect 43720 32564 43772 32570
rect 43720 32506 43772 32512
rect 43732 32434 43760 32506
rect 43720 32428 43772 32434
rect 43720 32370 43772 32376
rect 43732 31346 43760 32370
rect 43720 31340 43772 31346
rect 43720 31282 43772 31288
rect 43720 30660 43772 30666
rect 43720 30602 43772 30608
rect 43732 28218 43760 30602
rect 43824 29578 43852 34711
rect 43916 34202 43944 34886
rect 44100 34610 44128 35498
rect 44088 34604 44140 34610
rect 44088 34546 44140 34552
rect 44192 34490 44220 35634
rect 44008 34462 44220 34490
rect 43904 34196 43956 34202
rect 43904 34138 43956 34144
rect 43916 33522 43944 34138
rect 43904 33516 43956 33522
rect 43904 33458 43956 33464
rect 43904 32020 43956 32026
rect 43904 31962 43956 31968
rect 43916 30734 43944 31962
rect 43904 30728 43956 30734
rect 43904 30670 43956 30676
rect 43812 29572 43864 29578
rect 43812 29514 43864 29520
rect 43824 29102 43852 29514
rect 43916 29170 43944 30670
rect 44008 29646 44036 34462
rect 44180 34400 44232 34406
rect 44180 34342 44232 34348
rect 44192 34066 44220 34342
rect 44180 34060 44232 34066
rect 44180 34002 44232 34008
rect 44088 32904 44140 32910
rect 44088 32846 44140 32852
rect 44100 31346 44128 32846
rect 44284 31822 44312 35974
rect 44468 35834 44496 36110
rect 44928 36106 44956 36246
rect 45020 36242 45048 37062
rect 45192 36780 45244 36786
rect 45192 36722 45244 36728
rect 45100 36576 45152 36582
rect 45100 36518 45152 36524
rect 45008 36236 45060 36242
rect 45008 36178 45060 36184
rect 44916 36100 44968 36106
rect 44916 36042 44968 36048
rect 44456 35828 44508 35834
rect 44456 35770 44508 35776
rect 44456 34944 44508 34950
rect 44456 34886 44508 34892
rect 44468 34746 44496 34886
rect 44456 34740 44508 34746
rect 44456 34682 44508 34688
rect 45112 34542 45140 36518
rect 45204 36038 45232 36722
rect 45192 36032 45244 36038
rect 45192 35974 45244 35980
rect 45192 35692 45244 35698
rect 45192 35634 45244 35640
rect 45204 34950 45232 35634
rect 45192 34944 45244 34950
rect 45192 34886 45244 34892
rect 45100 34536 45152 34542
rect 45100 34478 45152 34484
rect 44548 34400 44600 34406
rect 44548 34342 44600 34348
rect 44560 33522 44588 34342
rect 44548 33516 44600 33522
rect 44548 33458 44600 33464
rect 44640 33516 44692 33522
rect 44640 33458 44692 33464
rect 44456 32768 44508 32774
rect 44456 32710 44508 32716
rect 44468 32502 44496 32710
rect 44456 32496 44508 32502
rect 44456 32438 44508 32444
rect 44272 31816 44324 31822
rect 44272 31758 44324 31764
rect 44088 31340 44140 31346
rect 44088 31282 44140 31288
rect 44100 29646 44128 31282
rect 44284 30938 44312 31758
rect 44560 31754 44588 33458
rect 44652 32978 44680 33458
rect 45204 33318 45232 34886
rect 45192 33312 45244 33318
rect 45192 33254 45244 33260
rect 44640 32972 44692 32978
rect 44640 32914 44692 32920
rect 44468 31726 44588 31754
rect 44272 30932 44324 30938
rect 44272 30874 44324 30880
rect 44180 30592 44232 30598
rect 44180 30534 44232 30540
rect 43996 29640 44048 29646
rect 43994 29608 43996 29617
rect 44088 29640 44140 29646
rect 44048 29608 44050 29617
rect 44088 29582 44140 29588
rect 43994 29543 44050 29552
rect 44100 29238 44128 29582
rect 44088 29232 44140 29238
rect 44088 29174 44140 29180
rect 43904 29164 43956 29170
rect 43904 29106 43956 29112
rect 43812 29096 43864 29102
rect 43812 29038 43864 29044
rect 43720 28212 43772 28218
rect 43720 28154 43772 28160
rect 43916 28064 43944 29106
rect 43996 28076 44048 28082
rect 43916 28036 43996 28064
rect 43996 28018 44048 28024
rect 43812 28008 43864 28014
rect 43812 27950 43864 27956
rect 43628 26784 43680 26790
rect 43628 26726 43680 26732
rect 43628 26308 43680 26314
rect 43628 26250 43680 26256
rect 43640 26042 43668 26250
rect 43628 26036 43680 26042
rect 43628 25978 43680 25984
rect 43824 25498 43852 27950
rect 44100 27554 44128 29174
rect 44192 28218 44220 30534
rect 44272 29708 44324 29714
rect 44272 29650 44324 29656
rect 44284 29209 44312 29650
rect 44270 29200 44326 29209
rect 44270 29135 44326 29144
rect 44284 29102 44312 29135
rect 44272 29096 44324 29102
rect 44272 29038 44324 29044
rect 44272 28416 44324 28422
rect 44272 28358 44324 28364
rect 44180 28212 44232 28218
rect 44180 28154 44232 28160
rect 44284 28082 44312 28358
rect 44272 28076 44324 28082
rect 44324 28036 44404 28064
rect 44272 28018 44324 28024
rect 44376 27674 44404 28036
rect 44364 27668 44416 27674
rect 44364 27610 44416 27616
rect 44008 27526 44128 27554
rect 43904 27328 43956 27334
rect 43904 27270 43956 27276
rect 43916 26314 43944 27270
rect 44008 27062 44036 27526
rect 44088 27464 44140 27470
rect 44088 27406 44140 27412
rect 43996 27056 44048 27062
rect 43996 26998 44048 27004
rect 43904 26308 43956 26314
rect 43904 26250 43956 26256
rect 44008 25906 44036 26998
rect 44100 26586 44128 27406
rect 44088 26580 44140 26586
rect 44088 26522 44140 26528
rect 43996 25900 44048 25906
rect 43996 25842 44048 25848
rect 44376 25702 44404 27610
rect 44468 26994 44496 31726
rect 44652 31278 44680 32914
rect 45296 32774 45324 37878
rect 45284 32768 45336 32774
rect 45284 32710 45336 32716
rect 45296 31686 45324 32710
rect 45284 31680 45336 31686
rect 45284 31622 45336 31628
rect 45388 31385 45416 43114
rect 45560 42696 45612 42702
rect 45560 42638 45612 42644
rect 45572 42362 45600 42638
rect 45560 42356 45612 42362
rect 45560 42298 45612 42304
rect 45468 40520 45520 40526
rect 45468 40462 45520 40468
rect 45480 39302 45508 40462
rect 45560 39364 45612 39370
rect 45560 39306 45612 39312
rect 45468 39296 45520 39302
rect 45468 39238 45520 39244
rect 45572 38350 45600 39306
rect 45744 38820 45796 38826
rect 45744 38762 45796 38768
rect 45652 38752 45704 38758
rect 45652 38694 45704 38700
rect 45560 38344 45612 38350
rect 45560 38286 45612 38292
rect 45664 38214 45692 38694
rect 45756 38418 45784 38762
rect 45744 38412 45796 38418
rect 45744 38354 45796 38360
rect 45652 38208 45704 38214
rect 45652 38150 45704 38156
rect 45468 37120 45520 37126
rect 45468 37062 45520 37068
rect 45480 36786 45508 37062
rect 45468 36780 45520 36786
rect 45468 36722 45520 36728
rect 45480 35494 45508 36722
rect 45744 36236 45796 36242
rect 45744 36178 45796 36184
rect 45756 35834 45784 36178
rect 45744 35828 45796 35834
rect 45744 35770 45796 35776
rect 45468 35488 45520 35494
rect 45468 35430 45520 35436
rect 45480 33590 45508 35430
rect 45848 34610 45876 47058
rect 46202 45928 46258 45937
rect 46202 45863 46204 45872
rect 46256 45863 46258 45872
rect 46204 45834 46256 45840
rect 46296 44192 46348 44198
rect 46296 44134 46348 44140
rect 46308 43450 46336 44134
rect 46492 43994 46520 47602
rect 47860 47456 47912 47462
rect 47860 47398 47912 47404
rect 47400 47184 47452 47190
rect 47400 47126 47452 47132
rect 47032 46096 47084 46102
rect 47032 46038 47084 46044
rect 47044 45558 47072 46038
rect 47124 45892 47176 45898
rect 47124 45834 47176 45840
rect 47032 45552 47084 45558
rect 47032 45494 47084 45500
rect 46940 44396 46992 44402
rect 46940 44338 46992 44344
rect 46480 43988 46532 43994
rect 46480 43930 46532 43936
rect 46296 43444 46348 43450
rect 46296 43386 46348 43392
rect 46308 43178 46336 43386
rect 46296 43172 46348 43178
rect 46296 43114 46348 43120
rect 46952 43110 46980 44338
rect 47044 44010 47072 45494
rect 47136 45082 47164 45834
rect 47124 45076 47176 45082
rect 47176 45036 47256 45064
rect 47124 45018 47176 45024
rect 47228 44470 47256 45036
rect 47216 44464 47268 44470
rect 47216 44406 47268 44412
rect 47308 44396 47360 44402
rect 47308 44338 47360 44344
rect 47216 44192 47268 44198
rect 47216 44134 47268 44140
rect 47044 43982 47164 44010
rect 47032 43920 47084 43926
rect 47032 43862 47084 43868
rect 47044 43654 47072 43862
rect 47136 43722 47164 43982
rect 47228 43722 47256 44134
rect 47124 43716 47176 43722
rect 47124 43658 47176 43664
rect 47216 43716 47268 43722
rect 47216 43658 47268 43664
rect 47032 43648 47084 43654
rect 47032 43590 47084 43596
rect 47032 43308 47084 43314
rect 47136 43296 47164 43658
rect 47320 43314 47348 44338
rect 47084 43268 47164 43296
rect 47032 43250 47084 43256
rect 46940 43104 46992 43110
rect 46940 43046 46992 43052
rect 46952 42378 46980 43046
rect 47136 42838 47164 43268
rect 47308 43308 47360 43314
rect 47308 43250 47360 43256
rect 47216 42900 47268 42906
rect 47216 42842 47268 42848
rect 47124 42832 47176 42838
rect 47124 42774 47176 42780
rect 46952 42350 47164 42378
rect 47228 42362 47256 42842
rect 46952 42226 46980 42350
rect 46940 42220 46992 42226
rect 46940 42162 46992 42168
rect 46664 41132 46716 41138
rect 46664 41074 46716 41080
rect 46676 40526 46704 41074
rect 46664 40520 46716 40526
rect 46664 40462 46716 40468
rect 46676 39914 46704 40462
rect 47032 40044 47084 40050
rect 47032 39986 47084 39992
rect 46664 39908 46716 39914
rect 46664 39850 46716 39856
rect 47044 39438 47072 39986
rect 46940 39432 46992 39438
rect 46940 39374 46992 39380
rect 47032 39432 47084 39438
rect 47032 39374 47084 39380
rect 46952 38350 46980 39374
rect 47136 39114 47164 42350
rect 47216 42356 47268 42362
rect 47216 42298 47268 42304
rect 47320 42226 47348 43250
rect 47308 42220 47360 42226
rect 47308 42162 47360 42168
rect 47216 39364 47268 39370
rect 47216 39306 47268 39312
rect 47044 39098 47164 39114
rect 47032 39092 47164 39098
rect 47084 39086 47164 39092
rect 47032 39034 47084 39040
rect 47136 38826 47164 39086
rect 47228 38894 47256 39306
rect 47216 38888 47268 38894
rect 47216 38830 47268 38836
rect 47124 38820 47176 38826
rect 47124 38762 47176 38768
rect 47216 38548 47268 38554
rect 47320 38536 47348 42162
rect 47412 41614 47440 47126
rect 47872 46578 47900 47398
rect 47860 46572 47912 46578
rect 47860 46514 47912 46520
rect 48688 46572 48740 46578
rect 48688 46514 48740 46520
rect 48964 46572 49016 46578
rect 48964 46514 49016 46520
rect 48044 46436 48096 46442
rect 48044 46378 48096 46384
rect 47952 45348 48004 45354
rect 47952 45290 48004 45296
rect 47964 44878 47992 45290
rect 47952 44872 48004 44878
rect 47952 44814 48004 44820
rect 47676 44736 47728 44742
rect 47676 44678 47728 44684
rect 47492 43784 47544 43790
rect 47492 43726 47544 43732
rect 47504 43450 47532 43726
rect 47688 43722 47716 44678
rect 47676 43716 47728 43722
rect 47676 43658 47728 43664
rect 47492 43444 47544 43450
rect 47492 43386 47544 43392
rect 47952 43444 48004 43450
rect 47952 43386 48004 43392
rect 47964 43178 47992 43386
rect 47952 43172 48004 43178
rect 47952 43114 48004 43120
rect 48056 42702 48084 46378
rect 48700 45966 48728 46514
rect 48780 46504 48832 46510
rect 48780 46446 48832 46452
rect 48504 45960 48556 45966
rect 48504 45902 48556 45908
rect 48688 45960 48740 45966
rect 48688 45902 48740 45908
rect 48516 45626 48544 45902
rect 48792 45665 48820 46446
rect 48778 45656 48834 45665
rect 48504 45620 48556 45626
rect 48778 45591 48834 45600
rect 48504 45562 48556 45568
rect 48412 45416 48464 45422
rect 48412 45358 48464 45364
rect 48424 44538 48452 45358
rect 48412 44532 48464 44538
rect 48412 44474 48464 44480
rect 48504 44532 48556 44538
rect 48504 44474 48556 44480
rect 48136 44192 48188 44198
rect 48136 44134 48188 44140
rect 48044 42696 48096 42702
rect 48044 42638 48096 42644
rect 48148 42294 48176 44134
rect 48228 43920 48280 43926
rect 48228 43862 48280 43868
rect 48240 43314 48268 43862
rect 48320 43648 48372 43654
rect 48320 43590 48372 43596
rect 48228 43308 48280 43314
rect 48228 43250 48280 43256
rect 48240 43110 48268 43250
rect 48228 43104 48280 43110
rect 48228 43046 48280 43052
rect 48332 42906 48360 43590
rect 48516 43450 48544 44474
rect 48976 44402 49004 46514
rect 49332 45824 49384 45830
rect 49332 45766 49384 45772
rect 49516 45824 49568 45830
rect 49516 45766 49568 45772
rect 50804 45824 50856 45830
rect 50804 45766 50856 45772
rect 52092 45824 52144 45830
rect 52092 45766 52144 45772
rect 49344 45354 49372 45766
rect 49424 45484 49476 45490
rect 49424 45426 49476 45432
rect 49332 45348 49384 45354
rect 49332 45290 49384 45296
rect 49148 44736 49200 44742
rect 49148 44678 49200 44684
rect 49240 44736 49292 44742
rect 49240 44678 49292 44684
rect 48872 44396 48924 44402
rect 48872 44338 48924 44344
rect 48964 44396 49016 44402
rect 48964 44338 49016 44344
rect 48780 43716 48832 43722
rect 48780 43658 48832 43664
rect 48504 43444 48556 43450
rect 48504 43386 48556 43392
rect 48596 43308 48648 43314
rect 48596 43250 48648 43256
rect 48320 42900 48372 42906
rect 48320 42842 48372 42848
rect 48412 42900 48464 42906
rect 48412 42842 48464 42848
rect 48228 42628 48280 42634
rect 48228 42570 48280 42576
rect 47860 42288 47912 42294
rect 47860 42230 47912 42236
rect 48136 42288 48188 42294
rect 48136 42230 48188 42236
rect 47492 42016 47544 42022
rect 47492 41958 47544 41964
rect 47504 41682 47532 41958
rect 47584 41812 47636 41818
rect 47584 41754 47636 41760
rect 47492 41676 47544 41682
rect 47492 41618 47544 41624
rect 47400 41608 47452 41614
rect 47400 41550 47452 41556
rect 47492 40384 47544 40390
rect 47492 40326 47544 40332
rect 47504 40186 47532 40326
rect 47492 40180 47544 40186
rect 47492 40122 47544 40128
rect 47596 39098 47624 41754
rect 47872 41274 47900 42230
rect 48044 42220 48096 42226
rect 48044 42162 48096 42168
rect 48056 42090 48084 42162
rect 48044 42084 48096 42090
rect 48044 42026 48096 42032
rect 48148 41818 48176 42230
rect 48240 42226 48268 42570
rect 48228 42220 48280 42226
rect 48228 42162 48280 42168
rect 48136 41812 48188 41818
rect 48136 41754 48188 41760
rect 48332 41614 48360 42842
rect 48424 42090 48452 42842
rect 48412 42084 48464 42090
rect 48412 42026 48464 42032
rect 48320 41608 48372 41614
rect 48320 41550 48372 41556
rect 47952 41472 48004 41478
rect 47952 41414 48004 41420
rect 47860 41268 47912 41274
rect 47860 41210 47912 41216
rect 47676 39840 47728 39846
rect 47676 39782 47728 39788
rect 47584 39092 47636 39098
rect 47584 39034 47636 39040
rect 47268 38508 47348 38536
rect 47688 38978 47716 39782
rect 47688 38950 47900 38978
rect 47216 38490 47268 38496
rect 47228 38418 47256 38490
rect 47216 38412 47268 38418
rect 47216 38354 47268 38360
rect 46940 38344 46992 38350
rect 46940 38286 46992 38292
rect 46952 37874 46980 38286
rect 47688 38214 47716 38950
rect 47872 38894 47900 38950
rect 47768 38888 47820 38894
rect 47768 38830 47820 38836
rect 47860 38888 47912 38894
rect 47860 38830 47912 38836
rect 47780 38282 47808 38830
rect 47860 38752 47912 38758
rect 47860 38694 47912 38700
rect 47964 38706 47992 41414
rect 48228 41268 48280 41274
rect 48228 41210 48280 41216
rect 48136 40656 48188 40662
rect 48136 40598 48188 40604
rect 48148 39302 48176 40598
rect 48240 40474 48268 41210
rect 48332 41138 48360 41550
rect 48320 41132 48372 41138
rect 48320 41074 48372 41080
rect 48332 40594 48360 41074
rect 48424 41002 48452 42026
rect 48608 41414 48636 43250
rect 48688 42764 48740 42770
rect 48688 42706 48740 42712
rect 48700 42294 48728 42706
rect 48688 42288 48740 42294
rect 48688 42230 48740 42236
rect 48792 41546 48820 43658
rect 48884 43178 48912 44338
rect 48964 44260 49016 44266
rect 48964 44202 49016 44208
rect 48976 43858 49004 44202
rect 49160 43858 49188 44678
rect 49252 44538 49280 44678
rect 49240 44532 49292 44538
rect 49240 44474 49292 44480
rect 49252 44402 49280 44474
rect 49240 44396 49292 44402
rect 49240 44338 49292 44344
rect 49240 44192 49292 44198
rect 49240 44134 49292 44140
rect 48964 43852 49016 43858
rect 48964 43794 49016 43800
rect 49148 43852 49200 43858
rect 49148 43794 49200 43800
rect 48872 43172 48924 43178
rect 48872 43114 48924 43120
rect 48976 43110 49004 43794
rect 49252 43790 49280 44134
rect 49240 43784 49292 43790
rect 49240 43726 49292 43732
rect 49344 43636 49372 45290
rect 49436 44946 49464 45426
rect 49424 44940 49476 44946
rect 49424 44882 49476 44888
rect 49160 43608 49372 43636
rect 48964 43104 49016 43110
rect 48964 43046 49016 43052
rect 48872 42900 48924 42906
rect 48872 42842 48924 42848
rect 48884 42702 48912 42842
rect 48872 42696 48924 42702
rect 48872 42638 48924 42644
rect 48976 42362 49004 43046
rect 48964 42356 49016 42362
rect 48964 42298 49016 42304
rect 49056 42356 49108 42362
rect 49056 42298 49108 42304
rect 48872 42288 48924 42294
rect 48872 42230 48924 42236
rect 48780 41540 48832 41546
rect 48780 41482 48832 41488
rect 48516 41386 48636 41414
rect 48412 40996 48464 41002
rect 48412 40938 48464 40944
rect 48412 40656 48464 40662
rect 48412 40598 48464 40604
rect 48320 40588 48372 40594
rect 48320 40530 48372 40536
rect 48424 40474 48452 40598
rect 48240 40446 48452 40474
rect 48320 40384 48372 40390
rect 48320 40326 48372 40332
rect 48332 40118 48360 40326
rect 48320 40112 48372 40118
rect 48320 40054 48372 40060
rect 48320 39976 48372 39982
rect 48318 39944 48320 39953
rect 48372 39944 48374 39953
rect 48318 39879 48374 39888
rect 48424 39370 48452 40446
rect 48516 39438 48544 41386
rect 48884 41070 48912 42230
rect 49068 42022 49096 42298
rect 49056 42016 49108 42022
rect 49056 41958 49108 41964
rect 49068 41818 49096 41958
rect 49056 41812 49108 41818
rect 49056 41754 49108 41760
rect 49056 41608 49108 41614
rect 49056 41550 49108 41556
rect 48872 41064 48924 41070
rect 48872 41006 48924 41012
rect 48964 40928 49016 40934
rect 48964 40870 49016 40876
rect 48976 40526 49004 40870
rect 48780 40520 48832 40526
rect 48780 40462 48832 40468
rect 48964 40520 49016 40526
rect 48964 40462 49016 40468
rect 48504 39432 48556 39438
rect 48504 39374 48556 39380
rect 48320 39364 48372 39370
rect 48320 39306 48372 39312
rect 48412 39364 48464 39370
rect 48412 39306 48464 39312
rect 48136 39296 48188 39302
rect 48136 39238 48188 39244
rect 48148 39030 48176 39238
rect 48332 39080 48360 39306
rect 48412 39092 48464 39098
rect 48332 39052 48412 39080
rect 48412 39034 48464 39040
rect 48136 39024 48188 39030
rect 48136 38966 48188 38972
rect 48320 38956 48372 38962
rect 48320 38898 48372 38904
rect 47768 38276 47820 38282
rect 47768 38218 47820 38224
rect 47676 38208 47728 38214
rect 47676 38150 47728 38156
rect 47780 37874 47808 38218
rect 46112 37868 46164 37874
rect 46112 37810 46164 37816
rect 46940 37868 46992 37874
rect 46940 37810 46992 37816
rect 47768 37868 47820 37874
rect 47768 37810 47820 37816
rect 46020 37800 46072 37806
rect 46020 37742 46072 37748
rect 46032 37262 46060 37742
rect 46124 37262 46152 37810
rect 46480 37664 46532 37670
rect 46480 37606 46532 37612
rect 46020 37256 46072 37262
rect 46020 37198 46072 37204
rect 46112 37256 46164 37262
rect 46112 37198 46164 37204
rect 46032 36786 46060 37198
rect 46020 36780 46072 36786
rect 46020 36722 46072 36728
rect 46124 36718 46152 37198
rect 46296 36780 46348 36786
rect 46296 36722 46348 36728
rect 46112 36712 46164 36718
rect 46112 36654 46164 36660
rect 46124 35766 46152 36654
rect 46308 36582 46336 36722
rect 46296 36576 46348 36582
rect 46296 36518 46348 36524
rect 46308 36088 46336 36518
rect 46492 36174 46520 37606
rect 46952 37466 46980 37810
rect 46940 37460 46992 37466
rect 46940 37402 46992 37408
rect 46952 37262 46980 37402
rect 46572 37256 46624 37262
rect 46572 37198 46624 37204
rect 46940 37256 46992 37262
rect 46940 37198 46992 37204
rect 46584 36786 46612 37198
rect 47780 37194 47808 37810
rect 47768 37188 47820 37194
rect 47768 37130 47820 37136
rect 47780 36854 47808 37130
rect 47872 37126 47900 38694
rect 47964 38678 48084 38706
rect 47860 37120 47912 37126
rect 47860 37062 47912 37068
rect 47768 36848 47820 36854
rect 47768 36790 47820 36796
rect 46572 36780 46624 36786
rect 46572 36722 46624 36728
rect 46480 36168 46532 36174
rect 46480 36110 46532 36116
rect 46216 36060 46336 36088
rect 46112 35760 46164 35766
rect 46112 35702 46164 35708
rect 46216 35698 46244 36060
rect 46584 36038 46612 36722
rect 46848 36712 46900 36718
rect 46848 36654 46900 36660
rect 46860 36174 46888 36654
rect 47400 36576 47452 36582
rect 47400 36518 47452 36524
rect 47584 36576 47636 36582
rect 47584 36518 47636 36524
rect 46940 36304 46992 36310
rect 46940 36246 46992 36252
rect 46848 36168 46900 36174
rect 46848 36110 46900 36116
rect 46572 36032 46624 36038
rect 46572 35974 46624 35980
rect 45928 35692 45980 35698
rect 45928 35634 45980 35640
rect 46204 35692 46256 35698
rect 46204 35634 46256 35640
rect 45940 35154 45968 35634
rect 46216 35562 46244 35634
rect 46204 35556 46256 35562
rect 46204 35498 46256 35504
rect 45928 35148 45980 35154
rect 45928 35090 45980 35096
rect 45940 34678 45968 35090
rect 45928 34672 45980 34678
rect 45928 34614 45980 34620
rect 45836 34604 45888 34610
rect 45836 34546 45888 34552
rect 45836 34196 45888 34202
rect 45836 34138 45888 34144
rect 45560 34128 45612 34134
rect 45560 34070 45612 34076
rect 45468 33584 45520 33590
rect 45468 33526 45520 33532
rect 45572 31754 45600 34070
rect 45848 33998 45876 34138
rect 45836 33992 45888 33998
rect 45836 33934 45888 33940
rect 45940 33318 45968 34614
rect 46584 34610 46612 35974
rect 46664 35488 46716 35494
rect 46664 35430 46716 35436
rect 46676 35086 46704 35430
rect 46952 35086 46980 36246
rect 47412 36174 47440 36518
rect 47596 36174 47624 36518
rect 47952 36304 48004 36310
rect 47952 36246 48004 36252
rect 47400 36168 47452 36174
rect 47400 36110 47452 36116
rect 47584 36168 47636 36174
rect 47584 36110 47636 36116
rect 47124 35624 47176 35630
rect 47124 35566 47176 35572
rect 47308 35624 47360 35630
rect 47308 35566 47360 35572
rect 46664 35080 46716 35086
rect 46664 35022 46716 35028
rect 46940 35080 46992 35086
rect 46940 35022 46992 35028
rect 46940 34944 46992 34950
rect 46992 34904 47072 34932
rect 46940 34886 46992 34892
rect 46112 34604 46164 34610
rect 46032 34564 46112 34592
rect 46032 33522 46060 34564
rect 46112 34546 46164 34552
rect 46572 34604 46624 34610
rect 46572 34546 46624 34552
rect 46296 34400 46348 34406
rect 46296 34342 46348 34348
rect 46204 33856 46256 33862
rect 46204 33798 46256 33804
rect 46020 33516 46072 33522
rect 46020 33458 46072 33464
rect 45928 33312 45980 33318
rect 45928 33254 45980 33260
rect 45940 32502 45968 33254
rect 45928 32496 45980 32502
rect 45928 32438 45980 32444
rect 46032 32366 46060 33458
rect 46216 32978 46244 33798
rect 46204 32972 46256 32978
rect 46204 32914 46256 32920
rect 46020 32360 46072 32366
rect 46020 32302 46072 32308
rect 45926 31920 45982 31929
rect 45926 31855 45982 31864
rect 45940 31822 45968 31855
rect 45928 31816 45980 31822
rect 45928 31758 45980 31764
rect 45560 31748 45612 31754
rect 45560 31690 45612 31696
rect 45940 31482 45968 31758
rect 46020 31748 46072 31754
rect 46020 31690 46072 31696
rect 45928 31476 45980 31482
rect 45928 31418 45980 31424
rect 46032 31414 46060 31690
rect 46020 31408 46072 31414
rect 45374 31376 45430 31385
rect 45192 31340 45244 31346
rect 46020 31350 46072 31356
rect 45374 31311 45430 31320
rect 45192 31282 45244 31288
rect 44640 31272 44692 31278
rect 44640 31214 44692 31220
rect 45204 30326 45232 31282
rect 45284 30660 45336 30666
rect 45284 30602 45336 30608
rect 45192 30320 45244 30326
rect 45192 30262 45244 30268
rect 44548 30252 44600 30258
rect 44548 30194 44600 30200
rect 44560 29850 44588 30194
rect 45296 30190 45324 30602
rect 45388 30376 45416 31311
rect 46204 31272 46256 31278
rect 46204 31214 46256 31220
rect 45928 30728 45980 30734
rect 45928 30670 45980 30676
rect 46112 30728 46164 30734
rect 46112 30670 46164 30676
rect 45388 30348 45600 30376
rect 45572 30258 45600 30348
rect 45744 30320 45796 30326
rect 45744 30262 45796 30268
rect 45560 30252 45612 30258
rect 45560 30194 45612 30200
rect 45284 30184 45336 30190
rect 45284 30126 45336 30132
rect 44548 29844 44600 29850
rect 44548 29786 44600 29792
rect 45192 29640 45244 29646
rect 45192 29582 45244 29588
rect 45284 29640 45336 29646
rect 45284 29582 45336 29588
rect 45098 29472 45154 29481
rect 45098 29407 45154 29416
rect 45112 29170 45140 29407
rect 45100 29164 45152 29170
rect 45100 29106 45152 29112
rect 44732 29028 44784 29034
rect 44732 28970 44784 28976
rect 44744 28694 44772 28970
rect 44732 28688 44784 28694
rect 44732 28630 44784 28636
rect 45008 28008 45060 28014
rect 45008 27950 45060 27956
rect 44824 27328 44876 27334
rect 44824 27270 44876 27276
rect 44836 26994 44864 27270
rect 44456 26988 44508 26994
rect 44456 26930 44508 26936
rect 44824 26988 44876 26994
rect 44824 26930 44876 26936
rect 45020 26382 45048 27950
rect 45112 27062 45140 29106
rect 45204 28762 45232 29582
rect 45296 28762 45324 29582
rect 45756 29578 45784 30262
rect 45468 29572 45520 29578
rect 45468 29514 45520 29520
rect 45744 29572 45796 29578
rect 45744 29514 45796 29520
rect 45480 29481 45508 29514
rect 45466 29472 45522 29481
rect 45466 29407 45522 29416
rect 45192 28756 45244 28762
rect 45192 28698 45244 28704
rect 45284 28756 45336 28762
rect 45284 28698 45336 28704
rect 45192 28620 45244 28626
rect 45192 28562 45244 28568
rect 45204 28490 45232 28562
rect 45192 28484 45244 28490
rect 45192 28426 45244 28432
rect 45296 28150 45324 28698
rect 45652 28552 45704 28558
rect 45652 28494 45704 28500
rect 45468 28212 45520 28218
rect 45468 28154 45520 28160
rect 45284 28144 45336 28150
rect 45284 28086 45336 28092
rect 45284 28008 45336 28014
rect 45284 27950 45336 27956
rect 45296 27674 45324 27950
rect 45376 27872 45428 27878
rect 45376 27814 45428 27820
rect 45284 27668 45336 27674
rect 45284 27610 45336 27616
rect 45388 27470 45416 27814
rect 45480 27470 45508 28154
rect 45664 28082 45692 28494
rect 45652 28076 45704 28082
rect 45652 28018 45704 28024
rect 45376 27464 45428 27470
rect 45376 27406 45428 27412
rect 45468 27464 45520 27470
rect 45468 27406 45520 27412
rect 45558 27296 45614 27305
rect 45558 27231 45614 27240
rect 45572 27130 45600 27231
rect 45560 27124 45612 27130
rect 45560 27066 45612 27072
rect 45664 27062 45692 28018
rect 45100 27056 45152 27062
rect 45100 26998 45152 27004
rect 45652 27056 45704 27062
rect 45652 26998 45704 27004
rect 45756 26994 45784 29514
rect 45834 29336 45890 29345
rect 45834 29271 45890 29280
rect 45848 28558 45876 29271
rect 45940 28937 45968 30670
rect 46020 30592 46072 30598
rect 46020 30534 46072 30540
rect 45926 28928 45982 28937
rect 45926 28863 45982 28872
rect 45836 28552 45888 28558
rect 45836 28494 45888 28500
rect 45744 26988 45796 26994
rect 45744 26930 45796 26936
rect 45848 26926 45876 28494
rect 45940 28014 45968 28863
rect 45928 28008 45980 28014
rect 45928 27950 45980 27956
rect 46032 27282 46060 30534
rect 46124 29714 46152 30670
rect 46112 29708 46164 29714
rect 46112 29650 46164 29656
rect 46124 29170 46152 29650
rect 46216 29238 46244 31214
rect 46308 30122 46336 34342
rect 46388 34060 46440 34066
rect 46388 34002 46440 34008
rect 46400 33386 46428 34002
rect 46388 33380 46440 33386
rect 46388 33322 46440 33328
rect 47044 33318 47072 34904
rect 47032 33312 47084 33318
rect 47032 33254 47084 33260
rect 46848 32904 46900 32910
rect 46848 32846 46900 32852
rect 46860 32434 46888 32846
rect 46940 32564 46992 32570
rect 46940 32506 46992 32512
rect 46848 32428 46900 32434
rect 46848 32370 46900 32376
rect 46952 32026 46980 32506
rect 46940 32020 46992 32026
rect 46940 31962 46992 31968
rect 46388 31680 46440 31686
rect 47044 31668 47072 33254
rect 47136 32366 47164 35566
rect 47320 35290 47348 35566
rect 47308 35284 47360 35290
rect 47308 35226 47360 35232
rect 47596 35018 47624 36110
rect 47964 36038 47992 36246
rect 47952 36032 48004 36038
rect 47952 35974 48004 35980
rect 47952 35692 48004 35698
rect 47952 35634 48004 35640
rect 47860 35148 47912 35154
rect 47860 35090 47912 35096
rect 47584 35012 47636 35018
rect 47584 34954 47636 34960
rect 47216 33652 47268 33658
rect 47216 33594 47268 33600
rect 47228 32570 47256 33594
rect 47398 33144 47454 33153
rect 47398 33079 47454 33088
rect 47412 32910 47440 33079
rect 47596 32978 47624 34954
rect 47872 34610 47900 35090
rect 47964 34950 47992 35634
rect 47952 34944 48004 34950
rect 47952 34886 48004 34892
rect 47860 34604 47912 34610
rect 47860 34546 47912 34552
rect 47860 34400 47912 34406
rect 47860 34342 47912 34348
rect 47768 33924 47820 33930
rect 47872 33912 47900 34342
rect 47820 33884 47900 33912
rect 47768 33866 47820 33872
rect 47872 33386 47900 33884
rect 47860 33380 47912 33386
rect 47860 33322 47912 33328
rect 47964 33266 47992 34886
rect 47872 33238 47992 33266
rect 47584 32972 47636 32978
rect 47584 32914 47636 32920
rect 47400 32904 47452 32910
rect 47400 32846 47452 32852
rect 47216 32564 47268 32570
rect 47216 32506 47268 32512
rect 47124 32360 47176 32366
rect 47124 32302 47176 32308
rect 47228 31890 47256 32506
rect 47596 31958 47624 32914
rect 47768 32020 47820 32026
rect 47768 31962 47820 31968
rect 47584 31952 47636 31958
rect 47584 31894 47636 31900
rect 47216 31884 47268 31890
rect 47216 31826 47268 31832
rect 47676 31884 47728 31890
rect 47676 31826 47728 31832
rect 47228 31754 47256 31826
rect 47228 31726 47348 31754
rect 47124 31680 47176 31686
rect 47044 31640 47124 31668
rect 46388 31622 46440 31628
rect 47124 31622 47176 31628
rect 46296 30116 46348 30122
rect 46296 30058 46348 30064
rect 46204 29232 46256 29238
rect 46204 29174 46256 29180
rect 46112 29164 46164 29170
rect 46112 29106 46164 29112
rect 46112 28416 46164 28422
rect 46112 28358 46164 28364
rect 46124 27470 46152 28358
rect 46112 27464 46164 27470
rect 46112 27406 46164 27412
rect 46032 27254 46152 27282
rect 45836 26920 45888 26926
rect 45836 26862 45888 26868
rect 45848 26586 45876 26862
rect 45836 26580 45888 26586
rect 45836 26522 45888 26528
rect 45008 26376 45060 26382
rect 45008 26318 45060 26324
rect 45928 26308 45980 26314
rect 45928 26250 45980 26256
rect 45836 26240 45888 26246
rect 45836 26182 45888 26188
rect 45848 25906 45876 26182
rect 45836 25900 45888 25906
rect 45836 25842 45888 25848
rect 45940 25838 45968 26250
rect 46020 25900 46072 25906
rect 46020 25842 46072 25848
rect 45928 25832 45980 25838
rect 45928 25774 45980 25780
rect 44180 25696 44232 25702
rect 44180 25638 44232 25644
rect 44364 25696 44416 25702
rect 44364 25638 44416 25644
rect 44916 25696 44968 25702
rect 44916 25638 44968 25644
rect 43812 25492 43864 25498
rect 43812 25434 43864 25440
rect 43168 25424 43220 25430
rect 43168 25366 43220 25372
rect 43076 25220 43128 25226
rect 43076 25162 43128 25168
rect 43088 24410 43116 25162
rect 44192 24750 44220 25638
rect 44180 24744 44232 24750
rect 44180 24686 44232 24692
rect 44928 24410 44956 25638
rect 45100 25288 45152 25294
rect 45100 25230 45152 25236
rect 43076 24404 43128 24410
rect 43076 24346 43128 24352
rect 44916 24404 44968 24410
rect 44916 24346 44968 24352
rect 45112 24206 45140 25230
rect 45192 25152 45244 25158
rect 45192 25094 45244 25100
rect 45204 24818 45232 25094
rect 45940 24886 45968 25774
rect 45928 24880 45980 24886
rect 45928 24822 45980 24828
rect 45192 24812 45244 24818
rect 45192 24754 45244 24760
rect 45376 24812 45428 24818
rect 45376 24754 45428 24760
rect 45388 24342 45416 24754
rect 45376 24336 45428 24342
rect 45376 24278 45428 24284
rect 43444 24200 43496 24206
rect 43444 24142 43496 24148
rect 45100 24200 45152 24206
rect 45100 24142 45152 24148
rect 43456 23730 43484 24142
rect 45284 24064 45336 24070
rect 45284 24006 45336 24012
rect 45296 23798 45324 24006
rect 46032 23798 46060 25842
rect 46124 24018 46152 27254
rect 46216 25294 46244 29174
rect 46308 29170 46336 30058
rect 46400 29850 46428 31622
rect 46848 31408 46900 31414
rect 46848 31350 46900 31356
rect 46938 31376 46994 31385
rect 46572 30932 46624 30938
rect 46572 30874 46624 30880
rect 46584 30734 46612 30874
rect 46572 30728 46624 30734
rect 46756 30728 46808 30734
rect 46572 30670 46624 30676
rect 46754 30696 46756 30705
rect 46808 30696 46810 30705
rect 46388 29844 46440 29850
rect 46388 29786 46440 29792
rect 46296 29164 46348 29170
rect 46296 29106 46348 29112
rect 46480 29096 46532 29102
rect 46480 29038 46532 29044
rect 46296 28552 46348 28558
rect 46296 28494 46348 28500
rect 46308 28218 46336 28494
rect 46296 28212 46348 28218
rect 46296 28154 46348 28160
rect 46492 28082 46520 29038
rect 46388 28076 46440 28082
rect 46388 28018 46440 28024
rect 46480 28076 46532 28082
rect 46480 28018 46532 28024
rect 46584 28064 46612 30670
rect 46754 30631 46810 30640
rect 46860 30598 46888 31350
rect 46938 31311 46940 31320
rect 46992 31311 46994 31320
rect 46940 31282 46992 31288
rect 46940 31136 46992 31142
rect 46940 31078 46992 31084
rect 47032 31136 47084 31142
rect 47032 31078 47084 31084
rect 46848 30592 46900 30598
rect 46848 30534 46900 30540
rect 46846 30424 46902 30433
rect 46846 30359 46902 30368
rect 46860 30258 46888 30359
rect 46664 30252 46716 30258
rect 46664 30194 46716 30200
rect 46848 30252 46900 30258
rect 46848 30194 46900 30200
rect 46676 29850 46704 30194
rect 46664 29844 46716 29850
rect 46664 29786 46716 29792
rect 46848 29708 46900 29714
rect 46848 29650 46900 29656
rect 46664 29640 46716 29646
rect 46664 29582 46716 29588
rect 46676 28558 46704 29582
rect 46860 29102 46888 29650
rect 46952 29170 46980 31078
rect 47044 30841 47072 31078
rect 47030 30832 47086 30841
rect 47030 30767 47086 30776
rect 47032 29708 47084 29714
rect 47032 29650 47084 29656
rect 46940 29164 46992 29170
rect 46940 29106 46992 29112
rect 46848 29096 46900 29102
rect 46848 29038 46900 29044
rect 46860 28626 46888 29038
rect 47044 28966 47072 29650
rect 47032 28960 47084 28966
rect 47136 28937 47164 31622
rect 47216 31204 47268 31210
rect 47216 31146 47268 31152
rect 47228 29850 47256 31146
rect 47216 29844 47268 29850
rect 47216 29786 47268 29792
rect 47216 29708 47268 29714
rect 47216 29650 47268 29656
rect 47228 29481 47256 29650
rect 47214 29472 47270 29481
rect 47214 29407 47270 29416
rect 47032 28902 47084 28908
rect 47122 28928 47178 28937
rect 47122 28863 47178 28872
rect 46848 28620 46900 28626
rect 46848 28562 46900 28568
rect 46664 28552 46716 28558
rect 46664 28494 46716 28500
rect 46756 28416 46808 28422
rect 46756 28358 46808 28364
rect 46664 28076 46716 28082
rect 46584 28036 46664 28064
rect 46400 27674 46428 28018
rect 46388 27668 46440 27674
rect 46388 27610 46440 27616
rect 46296 26988 46348 26994
rect 46296 26930 46348 26936
rect 46308 26042 46336 26930
rect 46584 26858 46612 28036
rect 46664 28018 46716 28024
rect 46768 27470 46796 28358
rect 46860 27606 46888 28562
rect 47136 28218 47164 28863
rect 47320 28694 47348 31726
rect 47584 31680 47636 31686
rect 47584 31622 47636 31628
rect 47596 30734 47624 31622
rect 47688 31414 47716 31826
rect 47676 31408 47728 31414
rect 47676 31350 47728 31356
rect 47584 30728 47636 30734
rect 47584 30670 47636 30676
rect 47584 30592 47636 30598
rect 47584 30534 47636 30540
rect 47676 30592 47728 30598
rect 47676 30534 47728 30540
rect 47596 30433 47624 30534
rect 47582 30424 47638 30433
rect 47688 30394 47716 30534
rect 47582 30359 47638 30368
rect 47676 30388 47728 30394
rect 47676 30330 47728 30336
rect 47676 30184 47728 30190
rect 47676 30126 47728 30132
rect 47688 29850 47716 30126
rect 47676 29844 47728 29850
rect 47676 29786 47728 29792
rect 47584 29776 47636 29782
rect 47584 29718 47636 29724
rect 47400 29640 47452 29646
rect 47400 29582 47452 29588
rect 47308 28688 47360 28694
rect 47308 28630 47360 28636
rect 47308 28484 47360 28490
rect 47308 28426 47360 28432
rect 47124 28212 47176 28218
rect 47124 28154 47176 28160
rect 47124 27872 47176 27878
rect 47124 27814 47176 27820
rect 47136 27674 47164 27814
rect 47124 27668 47176 27674
rect 47124 27610 47176 27616
rect 46848 27600 46900 27606
rect 46848 27542 46900 27548
rect 46756 27464 46808 27470
rect 46756 27406 46808 27412
rect 46664 27056 46716 27062
rect 46664 26998 46716 27004
rect 46388 26852 46440 26858
rect 46388 26794 46440 26800
rect 46572 26852 46624 26858
rect 46572 26794 46624 26800
rect 46400 26246 46428 26794
rect 46676 26625 46704 26998
rect 46848 26988 46900 26994
rect 46848 26930 46900 26936
rect 46756 26920 46808 26926
rect 46756 26862 46808 26868
rect 46662 26616 46718 26625
rect 46662 26551 46718 26560
rect 46768 26450 46796 26862
rect 46860 26586 46888 26930
rect 47032 26784 47084 26790
rect 47032 26726 47084 26732
rect 46848 26580 46900 26586
rect 46848 26522 46900 26528
rect 46480 26444 46532 26450
rect 46480 26386 46532 26392
rect 46756 26444 46808 26450
rect 46756 26386 46808 26392
rect 46388 26240 46440 26246
rect 46388 26182 46440 26188
rect 46296 26036 46348 26042
rect 46296 25978 46348 25984
rect 46308 25498 46336 25978
rect 46296 25492 46348 25498
rect 46296 25434 46348 25440
rect 46204 25288 46256 25294
rect 46204 25230 46256 25236
rect 46216 24138 46244 25230
rect 46296 25152 46348 25158
rect 46296 25094 46348 25100
rect 46308 24274 46336 25094
rect 46296 24268 46348 24274
rect 46296 24210 46348 24216
rect 46204 24132 46256 24138
rect 46204 24074 46256 24080
rect 46296 24064 46348 24070
rect 46124 23990 46244 24018
rect 46296 24006 46348 24012
rect 45284 23792 45336 23798
rect 45284 23734 45336 23740
rect 46020 23792 46072 23798
rect 46020 23734 46072 23740
rect 43444 23724 43496 23730
rect 43444 23666 43496 23672
rect 42984 23520 43036 23526
rect 42984 23462 43036 23468
rect 42996 23118 43024 23462
rect 42984 23112 43036 23118
rect 42984 23054 43036 23060
rect 43456 23050 43484 23666
rect 46216 23050 46244 23990
rect 46308 23866 46336 24006
rect 46400 23866 46428 26182
rect 46492 25430 46520 26386
rect 46938 26072 46994 26081
rect 46938 26007 46940 26016
rect 46992 26007 46994 26016
rect 46940 25978 46992 25984
rect 47044 25906 47072 26726
rect 47136 26382 47164 27610
rect 47320 27334 47348 28426
rect 47412 28370 47440 29582
rect 47492 29164 47544 29170
rect 47492 29106 47544 29112
rect 47504 28558 47532 29106
rect 47492 28552 47544 28558
rect 47492 28494 47544 28500
rect 47412 28342 47532 28370
rect 47504 27334 47532 28342
rect 47308 27328 47360 27334
rect 47308 27270 47360 27276
rect 47492 27328 47544 27334
rect 47492 27270 47544 27276
rect 47216 26512 47268 26518
rect 47216 26454 47268 26460
rect 47124 26376 47176 26382
rect 47124 26318 47176 26324
rect 47136 25974 47164 26318
rect 47124 25968 47176 25974
rect 47124 25910 47176 25916
rect 47032 25900 47084 25906
rect 47032 25842 47084 25848
rect 46480 25424 46532 25430
rect 46480 25366 46532 25372
rect 47228 25294 47256 26454
rect 47504 26382 47532 27270
rect 47492 26376 47544 26382
rect 47492 26318 47544 26324
rect 47596 25974 47624 29718
rect 47676 29232 47728 29238
rect 47676 29174 47728 29180
rect 47688 28762 47716 29174
rect 47676 28756 47728 28762
rect 47676 28698 47728 28704
rect 47676 28552 47728 28558
rect 47676 28494 47728 28500
rect 47688 27674 47716 28494
rect 47676 27668 47728 27674
rect 47676 27610 47728 27616
rect 47676 26988 47728 26994
rect 47676 26930 47728 26936
rect 47688 26518 47716 26930
rect 47676 26512 47728 26518
rect 47676 26454 47728 26460
rect 47676 26308 47728 26314
rect 47676 26250 47728 26256
rect 47584 25968 47636 25974
rect 47584 25910 47636 25916
rect 47308 25492 47360 25498
rect 47308 25434 47360 25440
rect 47320 25294 47348 25434
rect 47032 25288 47084 25294
rect 47032 25230 47084 25236
rect 47216 25288 47268 25294
rect 47216 25230 47268 25236
rect 47308 25288 47360 25294
rect 47308 25230 47360 25236
rect 46940 25220 46992 25226
rect 46940 25162 46992 25168
rect 46952 24818 46980 25162
rect 46940 24812 46992 24818
rect 46940 24754 46992 24760
rect 46296 23860 46348 23866
rect 46296 23802 46348 23808
rect 46388 23860 46440 23866
rect 46388 23802 46440 23808
rect 46952 23730 46980 24754
rect 47044 24682 47072 25230
rect 47584 25152 47636 25158
rect 47584 25094 47636 25100
rect 47032 24676 47084 24682
rect 47032 24618 47084 24624
rect 47044 24410 47072 24618
rect 47596 24614 47624 25094
rect 47584 24608 47636 24614
rect 47584 24550 47636 24556
rect 47032 24404 47084 24410
rect 47032 24346 47084 24352
rect 47688 24274 47716 26250
rect 47676 24268 47728 24274
rect 47676 24210 47728 24216
rect 47400 24200 47452 24206
rect 47400 24142 47452 24148
rect 46940 23724 46992 23730
rect 46940 23666 46992 23672
rect 46848 23520 46900 23526
rect 46848 23462 46900 23468
rect 42800 23044 42852 23050
rect 42800 22986 42852 22992
rect 43444 23044 43496 23050
rect 43444 22986 43496 22992
rect 46204 23044 46256 23050
rect 46204 22986 46256 22992
rect 46480 23044 46532 23050
rect 46480 22986 46532 22992
rect 42812 22710 42840 22986
rect 43904 22976 43956 22982
rect 43904 22918 43956 22924
rect 44456 22976 44508 22982
rect 44456 22918 44508 22924
rect 43916 22778 43944 22918
rect 43904 22772 43956 22778
rect 43904 22714 43956 22720
rect 44468 22710 44496 22918
rect 46216 22710 46244 22986
rect 46492 22778 46520 22986
rect 46480 22772 46532 22778
rect 46480 22714 46532 22720
rect 42800 22704 42852 22710
rect 42800 22646 42852 22652
rect 44456 22704 44508 22710
rect 44456 22646 44508 22652
rect 46204 22704 46256 22710
rect 46204 22646 46256 22652
rect 46860 22642 46888 23462
rect 46952 23322 46980 23666
rect 47032 23588 47084 23594
rect 47032 23530 47084 23536
rect 46940 23316 46992 23322
rect 46940 23258 46992 23264
rect 42708 22636 42760 22642
rect 42708 22578 42760 22584
rect 46848 22636 46900 22642
rect 46848 22578 46900 22584
rect 39212 22092 39264 22098
rect 39212 22034 39264 22040
rect 47044 22030 47072 23530
rect 47412 23202 47440 24142
rect 47780 23730 47808 31962
rect 47872 31754 47900 33238
rect 47952 32768 48004 32774
rect 47952 32710 48004 32716
rect 47860 31748 47912 31754
rect 47860 31690 47912 31696
rect 47872 30734 47900 31690
rect 47860 30728 47912 30734
rect 47860 30670 47912 30676
rect 47964 29646 47992 32710
rect 48056 30818 48084 38678
rect 48332 38554 48360 38898
rect 48320 38548 48372 38554
rect 48320 38490 48372 38496
rect 48226 38040 48282 38049
rect 48226 37975 48282 37984
rect 48240 37874 48268 37975
rect 48320 37936 48372 37942
rect 48320 37878 48372 37884
rect 48228 37868 48280 37874
rect 48228 37810 48280 37816
rect 48332 37262 48360 37878
rect 48424 37874 48452 39034
rect 48516 37890 48544 39374
rect 48688 39296 48740 39302
rect 48688 39238 48740 39244
rect 48700 38214 48728 39238
rect 48688 38208 48740 38214
rect 48688 38150 48740 38156
rect 48700 37942 48728 38150
rect 48688 37936 48740 37942
rect 48516 37874 48636 37890
rect 48688 37878 48740 37884
rect 48412 37868 48464 37874
rect 48516 37868 48648 37874
rect 48516 37862 48596 37868
rect 48412 37810 48464 37816
rect 48596 37810 48648 37816
rect 48320 37256 48372 37262
rect 48320 37198 48372 37204
rect 48424 37194 48452 37810
rect 48608 37330 48636 37810
rect 48596 37324 48648 37330
rect 48596 37266 48648 37272
rect 48412 37188 48464 37194
rect 48412 37130 48464 37136
rect 48136 36644 48188 36650
rect 48136 36586 48188 36592
rect 48148 36038 48176 36586
rect 48424 36106 48452 37130
rect 48608 36922 48636 37266
rect 48688 37120 48740 37126
rect 48688 37062 48740 37068
rect 48596 36916 48648 36922
rect 48596 36858 48648 36864
rect 48700 36242 48728 37062
rect 48688 36236 48740 36242
rect 48688 36178 48740 36184
rect 48412 36100 48464 36106
rect 48412 36042 48464 36048
rect 48136 36032 48188 36038
rect 48136 35974 48188 35980
rect 48504 36032 48556 36038
rect 48504 35974 48556 35980
rect 48148 35086 48176 35974
rect 48320 35556 48372 35562
rect 48320 35498 48372 35504
rect 48332 35154 48360 35498
rect 48320 35148 48372 35154
rect 48320 35090 48372 35096
rect 48136 35080 48188 35086
rect 48136 35022 48188 35028
rect 48320 35012 48372 35018
rect 48320 34954 48372 34960
rect 48332 34610 48360 34954
rect 48320 34604 48372 34610
rect 48320 34546 48372 34552
rect 48332 33862 48360 34546
rect 48320 33856 48372 33862
rect 48320 33798 48372 33804
rect 48228 33516 48280 33522
rect 48228 33458 48280 33464
rect 48136 32224 48188 32230
rect 48136 32166 48188 32172
rect 48148 32026 48176 32166
rect 48136 32020 48188 32026
rect 48136 31962 48188 31968
rect 48240 31822 48268 33458
rect 48228 31816 48280 31822
rect 48228 31758 48280 31764
rect 48332 31482 48360 33798
rect 48516 33522 48544 35974
rect 48792 35850 48820 40462
rect 49068 40372 49096 41550
rect 49160 41449 49188 43608
rect 49424 42696 49476 42702
rect 49330 42664 49386 42673
rect 49424 42638 49476 42644
rect 49330 42599 49332 42608
rect 49384 42599 49386 42608
rect 49332 42570 49384 42576
rect 49240 42560 49292 42566
rect 49238 42528 49240 42537
rect 49292 42528 49294 42537
rect 49238 42463 49294 42472
rect 49240 42220 49292 42226
rect 49240 42162 49292 42168
rect 49252 41818 49280 42162
rect 49436 42090 49464 42638
rect 49424 42084 49476 42090
rect 49424 42026 49476 42032
rect 49240 41812 49292 41818
rect 49240 41754 49292 41760
rect 49240 41540 49292 41546
rect 49240 41482 49292 41488
rect 49146 41440 49202 41449
rect 49146 41375 49202 41384
rect 49252 41274 49280 41482
rect 49240 41268 49292 41274
rect 49240 41210 49292 41216
rect 49332 41132 49384 41138
rect 49332 41074 49384 41080
rect 48976 40344 49096 40372
rect 48872 39432 48924 39438
rect 48872 39374 48924 39380
rect 48884 39098 48912 39374
rect 48872 39092 48924 39098
rect 48872 39034 48924 39040
rect 48608 35822 48820 35850
rect 48608 34202 48636 35822
rect 48780 35692 48832 35698
rect 48780 35634 48832 35640
rect 48688 35556 48740 35562
rect 48688 35498 48740 35504
rect 48700 35086 48728 35498
rect 48688 35080 48740 35086
rect 48688 35022 48740 35028
rect 48700 34728 48728 35022
rect 48792 35018 48820 35634
rect 48872 35624 48924 35630
rect 48872 35566 48924 35572
rect 48884 35086 48912 35566
rect 48872 35080 48924 35086
rect 48872 35022 48924 35028
rect 48780 35012 48832 35018
rect 48780 34954 48832 34960
rect 48700 34700 48820 34728
rect 48688 34604 48740 34610
rect 48688 34546 48740 34552
rect 48596 34196 48648 34202
rect 48596 34138 48648 34144
rect 48700 33998 48728 34546
rect 48792 33998 48820 34700
rect 48884 34678 48912 35022
rect 48976 34746 49004 40344
rect 49344 39930 49372 41074
rect 49436 40458 49464 42026
rect 49528 40526 49556 45766
rect 50816 45354 50844 45766
rect 50896 45416 50948 45422
rect 50896 45358 50948 45364
rect 51540 45416 51592 45422
rect 51540 45358 51592 45364
rect 50804 45348 50856 45354
rect 50804 45290 50856 45296
rect 50528 45280 50580 45286
rect 50528 45222 50580 45228
rect 50540 44878 50568 45222
rect 50620 44940 50672 44946
rect 50620 44882 50672 44888
rect 50528 44872 50580 44878
rect 50528 44814 50580 44820
rect 50528 44736 50580 44742
rect 50528 44678 50580 44684
rect 50436 44396 50488 44402
rect 50436 44338 50488 44344
rect 50344 44192 50396 44198
rect 50344 44134 50396 44140
rect 49608 43852 49660 43858
rect 49608 43794 49660 43800
rect 49620 43314 49648 43794
rect 50356 43790 50384 44134
rect 50448 43994 50476 44338
rect 50540 44198 50568 44678
rect 50528 44192 50580 44198
rect 50528 44134 50580 44140
rect 50436 43988 50488 43994
rect 50436 43930 50488 43936
rect 50344 43784 50396 43790
rect 50344 43726 50396 43732
rect 50068 43648 50120 43654
rect 50448 43636 50476 43930
rect 50540 43790 50568 44134
rect 50632 43994 50660 44882
rect 50816 44266 50844 45290
rect 50908 45082 50936 45358
rect 50896 45076 50948 45082
rect 50896 45018 50948 45024
rect 51172 44464 51224 44470
rect 51172 44406 51224 44412
rect 50988 44328 51040 44334
rect 50988 44270 51040 44276
rect 50804 44260 50856 44266
rect 50804 44202 50856 44208
rect 50620 43988 50672 43994
rect 50620 43930 50672 43936
rect 50816 43926 50844 44202
rect 50804 43920 50856 43926
rect 50724 43880 50804 43908
rect 50528 43784 50580 43790
rect 50528 43726 50580 43732
rect 50724 43722 50752 43880
rect 50804 43862 50856 43868
rect 51000 43790 51028 44270
rect 50988 43784 51040 43790
rect 50988 43726 51040 43732
rect 50712 43716 50764 43722
rect 50632 43676 50712 43704
rect 50632 43636 50660 43676
rect 50712 43658 50764 43664
rect 50448 43608 50660 43636
rect 50896 43648 50948 43654
rect 50068 43590 50120 43596
rect 51184 43602 51212 44406
rect 51552 43858 51580 45358
rect 52000 44940 52052 44946
rect 52000 44882 52052 44888
rect 51724 44396 51776 44402
rect 51724 44338 51776 44344
rect 51632 44328 51684 44334
rect 51632 44270 51684 44276
rect 51540 43852 51592 43858
rect 51540 43794 51592 43800
rect 50948 43596 51212 43602
rect 50896 43590 51212 43596
rect 50080 43314 50108 43590
rect 50908 43574 51212 43590
rect 51552 43314 51580 43794
rect 51644 43772 51672 44270
rect 51736 43994 51764 44338
rect 51724 43988 51776 43994
rect 51724 43930 51776 43936
rect 51816 43784 51868 43790
rect 51644 43744 51816 43772
rect 51816 43726 51868 43732
rect 49608 43308 49660 43314
rect 49608 43250 49660 43256
rect 50068 43308 50120 43314
rect 50068 43250 50120 43256
rect 50528 43308 50580 43314
rect 50528 43250 50580 43256
rect 51540 43308 51592 43314
rect 51540 43250 51592 43256
rect 49976 43240 50028 43246
rect 49976 43182 50028 43188
rect 49988 42906 50016 43182
rect 49976 42900 50028 42906
rect 49976 42842 50028 42848
rect 49608 42832 49660 42838
rect 49608 42774 49660 42780
rect 49620 42226 49648 42774
rect 49884 42696 49936 42702
rect 49884 42638 49936 42644
rect 50342 42664 50398 42673
rect 49608 42220 49660 42226
rect 49608 42162 49660 42168
rect 49620 41546 49648 42162
rect 49700 42016 49752 42022
rect 49700 41958 49752 41964
rect 49712 41682 49740 41958
rect 49700 41676 49752 41682
rect 49700 41618 49752 41624
rect 49608 41540 49660 41546
rect 49608 41482 49660 41488
rect 49792 41472 49844 41478
rect 49606 41440 49662 41449
rect 49792 41414 49844 41420
rect 49606 41375 49662 41384
rect 49620 41138 49648 41375
rect 49608 41132 49660 41138
rect 49608 41074 49660 41080
rect 49608 40996 49660 41002
rect 49608 40938 49660 40944
rect 49516 40520 49568 40526
rect 49516 40462 49568 40468
rect 49424 40452 49476 40458
rect 49424 40394 49476 40400
rect 49528 40118 49556 40462
rect 49516 40112 49568 40118
rect 49516 40054 49568 40060
rect 49344 39902 49556 39930
rect 49620 39914 49648 40938
rect 49700 40384 49752 40390
rect 49700 40326 49752 40332
rect 49332 39296 49384 39302
rect 49332 39238 49384 39244
rect 49056 38956 49108 38962
rect 49056 38898 49108 38904
rect 49068 38418 49096 38898
rect 49344 38758 49372 39238
rect 49332 38752 49384 38758
rect 49332 38694 49384 38700
rect 49056 38412 49108 38418
rect 49056 38354 49108 38360
rect 49240 38412 49292 38418
rect 49240 38354 49292 38360
rect 49148 37120 49200 37126
rect 49148 37062 49200 37068
rect 49160 36718 49188 37062
rect 49252 36786 49280 38354
rect 49344 38049 49372 38694
rect 49424 38344 49476 38350
rect 49424 38286 49476 38292
rect 49330 38040 49386 38049
rect 49330 37975 49386 37984
rect 49332 37936 49384 37942
rect 49332 37878 49384 37884
rect 49344 37398 49372 37878
rect 49332 37392 49384 37398
rect 49332 37334 49384 37340
rect 49332 37256 49384 37262
rect 49332 37198 49384 37204
rect 49240 36780 49292 36786
rect 49240 36722 49292 36728
rect 49148 36712 49200 36718
rect 49148 36654 49200 36660
rect 49252 36378 49280 36722
rect 49240 36372 49292 36378
rect 49240 36314 49292 36320
rect 49056 36168 49108 36174
rect 49056 36110 49108 36116
rect 49068 35222 49096 36110
rect 49344 36038 49372 37198
rect 49332 36032 49384 36038
rect 49332 35974 49384 35980
rect 49056 35216 49108 35222
rect 49056 35158 49108 35164
rect 48964 34740 49016 34746
rect 48964 34682 49016 34688
rect 48872 34672 48924 34678
rect 48872 34614 48924 34620
rect 49332 34604 49384 34610
rect 49332 34546 49384 34552
rect 48688 33992 48740 33998
rect 48688 33934 48740 33940
rect 48780 33992 48832 33998
rect 48780 33934 48832 33940
rect 48596 33924 48648 33930
rect 48596 33866 48648 33872
rect 48504 33516 48556 33522
rect 48504 33458 48556 33464
rect 48412 33448 48464 33454
rect 48412 33390 48464 33396
rect 48424 33114 48452 33390
rect 48412 33108 48464 33114
rect 48412 33050 48464 33056
rect 48608 32910 48636 33866
rect 48688 33516 48740 33522
rect 48688 33458 48740 33464
rect 48596 32904 48648 32910
rect 48596 32846 48648 32852
rect 48412 32836 48464 32842
rect 48412 32778 48464 32784
rect 48424 32502 48452 32778
rect 48596 32768 48648 32774
rect 48596 32710 48648 32716
rect 48412 32496 48464 32502
rect 48412 32438 48464 32444
rect 48608 32434 48636 32710
rect 48596 32428 48648 32434
rect 48596 32370 48648 32376
rect 48608 31822 48636 32370
rect 48700 32026 48728 33458
rect 48792 33046 48820 33934
rect 49344 33930 49372 34546
rect 49332 33924 49384 33930
rect 49332 33866 49384 33872
rect 48780 33040 48832 33046
rect 48780 32982 48832 32988
rect 49436 32502 49464 38286
rect 49424 32496 49476 32502
rect 49424 32438 49476 32444
rect 49528 32230 49556 39902
rect 49608 39908 49660 39914
rect 49608 39850 49660 39856
rect 49712 39506 49740 40326
rect 49804 39574 49832 41414
rect 49896 40458 49924 42638
rect 50342 42599 50344 42608
rect 50396 42599 50398 42608
rect 50344 42570 50396 42576
rect 49976 42220 50028 42226
rect 49976 42162 50028 42168
rect 49988 41478 50016 42162
rect 50540 41614 50568 43250
rect 51448 43240 51500 43246
rect 51448 43182 51500 43188
rect 51264 42764 51316 42770
rect 51264 42706 51316 42712
rect 51276 42158 51304 42706
rect 51080 42152 51132 42158
rect 51080 42094 51132 42100
rect 51264 42152 51316 42158
rect 51264 42094 51316 42100
rect 51092 41818 51120 42094
rect 51080 41812 51132 41818
rect 51080 41754 51132 41760
rect 50528 41608 50580 41614
rect 50528 41550 50580 41556
rect 49976 41472 50028 41478
rect 49976 41414 50028 41420
rect 50896 41472 50948 41478
rect 50896 41414 50948 41420
rect 50988 41472 51040 41478
rect 50988 41414 51040 41420
rect 50252 41268 50304 41274
rect 50252 41210 50304 41216
rect 50264 41070 50292 41210
rect 50804 41132 50856 41138
rect 50804 41074 50856 41080
rect 50252 41064 50304 41070
rect 50252 41006 50304 41012
rect 49884 40452 49936 40458
rect 49884 40394 49936 40400
rect 50264 40050 50292 41006
rect 50252 40044 50304 40050
rect 50252 39986 50304 39992
rect 50160 39908 50212 39914
rect 50160 39850 50212 39856
rect 49792 39568 49844 39574
rect 49792 39510 49844 39516
rect 49700 39500 49752 39506
rect 49700 39442 49752 39448
rect 49974 38448 50030 38457
rect 49974 38383 50030 38392
rect 49792 37664 49844 37670
rect 49792 37606 49844 37612
rect 49700 37256 49752 37262
rect 49700 37198 49752 37204
rect 49712 36718 49740 37198
rect 49700 36712 49752 36718
rect 49700 36654 49752 36660
rect 49804 36258 49832 37606
rect 49988 36854 50016 38383
rect 50068 36916 50120 36922
rect 50068 36858 50120 36864
rect 49976 36848 50028 36854
rect 49976 36790 50028 36796
rect 50080 36582 50108 36858
rect 50068 36576 50120 36582
rect 50068 36518 50120 36524
rect 49712 36242 49832 36258
rect 49700 36236 49832 36242
rect 49752 36230 49832 36236
rect 49700 36178 49752 36184
rect 49712 35290 49740 36178
rect 50080 36106 50108 36518
rect 50068 36100 50120 36106
rect 50068 36042 50120 36048
rect 49976 35556 50028 35562
rect 49976 35498 50028 35504
rect 49700 35284 49752 35290
rect 49700 35226 49752 35232
rect 49988 35018 50016 35498
rect 49976 35012 50028 35018
rect 49976 34954 50028 34960
rect 49608 34672 49660 34678
rect 49608 34614 49660 34620
rect 49620 33998 49648 34614
rect 49976 34400 50028 34406
rect 49976 34342 50028 34348
rect 49988 34066 50016 34342
rect 49976 34060 50028 34066
rect 49976 34002 50028 34008
rect 49608 33992 49660 33998
rect 49608 33934 49660 33940
rect 49700 33924 49752 33930
rect 49700 33866 49752 33872
rect 49712 33658 49740 33866
rect 49700 33652 49752 33658
rect 49700 33594 49752 33600
rect 49988 33522 50016 34002
rect 49976 33516 50028 33522
rect 49976 33458 50028 33464
rect 49792 33448 49844 33454
rect 49792 33390 49844 33396
rect 49608 33312 49660 33318
rect 49608 33254 49660 33260
rect 49700 33312 49752 33318
rect 49700 33254 49752 33260
rect 49620 32910 49648 33254
rect 49608 32904 49660 32910
rect 49608 32846 49660 32852
rect 49516 32224 49568 32230
rect 49516 32166 49568 32172
rect 48688 32020 48740 32026
rect 48688 31962 48740 31968
rect 49056 32020 49108 32026
rect 49056 31962 49108 31968
rect 48596 31816 48648 31822
rect 48596 31758 48648 31764
rect 48320 31476 48372 31482
rect 48320 31418 48372 31424
rect 48320 31340 48372 31346
rect 48320 31282 48372 31288
rect 48056 30790 48268 30818
rect 48044 30728 48096 30734
rect 48044 30670 48096 30676
rect 48134 30696 48190 30705
rect 47952 29640 48004 29646
rect 47952 29582 48004 29588
rect 47860 29572 47912 29578
rect 47860 29514 47912 29520
rect 47872 29345 47900 29514
rect 47858 29336 47914 29345
rect 47858 29271 47914 29280
rect 47950 29200 48006 29209
rect 47950 29135 47952 29144
rect 48004 29135 48006 29144
rect 47952 29106 48004 29112
rect 47860 29028 47912 29034
rect 47860 28970 47912 28976
rect 47872 28422 47900 28970
rect 47860 28416 47912 28422
rect 47860 28358 47912 28364
rect 48056 28082 48084 30670
rect 48134 30631 48136 30640
rect 48188 30631 48190 30640
rect 48136 30602 48188 30608
rect 48136 29640 48188 29646
rect 48136 29582 48188 29588
rect 48148 29034 48176 29582
rect 48240 29209 48268 30790
rect 48332 30394 48360 31282
rect 48412 31204 48464 31210
rect 48412 31146 48464 31152
rect 48424 30802 48452 31146
rect 48412 30796 48464 30802
rect 48412 30738 48464 30744
rect 48320 30388 48372 30394
rect 48320 30330 48372 30336
rect 48608 30274 48636 31758
rect 48964 31272 49016 31278
rect 48964 31214 49016 31220
rect 48332 30258 48636 30274
rect 48976 30274 49004 31214
rect 49068 30734 49096 31962
rect 49608 31136 49660 31142
rect 49608 31078 49660 31084
rect 49056 30728 49108 30734
rect 49056 30670 49108 30676
rect 49620 30308 49648 31078
rect 49712 30666 49740 33254
rect 49804 33114 49832 33390
rect 49988 33318 50016 33458
rect 50068 33380 50120 33386
rect 50068 33322 50120 33328
rect 49976 33312 50028 33318
rect 49976 33254 50028 33260
rect 49792 33108 49844 33114
rect 49792 33050 49844 33056
rect 49792 32904 49844 32910
rect 49792 32846 49844 32852
rect 49804 32570 49832 32846
rect 49792 32564 49844 32570
rect 49792 32506 49844 32512
rect 49988 31754 50016 33254
rect 50080 33114 50108 33322
rect 50068 33108 50120 33114
rect 50068 33050 50120 33056
rect 49896 31726 50016 31754
rect 49896 31142 49924 31726
rect 49884 31136 49936 31142
rect 49884 31078 49936 31084
rect 49700 30660 49752 30666
rect 49700 30602 49752 30608
rect 49700 30320 49752 30326
rect 49620 30280 49700 30308
rect 48320 30252 48636 30258
rect 48372 30246 48636 30252
rect 48872 30252 48924 30258
rect 48320 30194 48372 30200
rect 48516 30190 48544 30246
rect 48976 30246 49188 30274
rect 49700 30262 49752 30268
rect 48872 30194 48924 30200
rect 48504 30184 48556 30190
rect 48504 30126 48556 30132
rect 48516 29646 48544 30126
rect 48504 29640 48556 29646
rect 48504 29582 48556 29588
rect 48320 29572 48372 29578
rect 48320 29514 48372 29520
rect 48226 29200 48282 29209
rect 48332 29170 48360 29514
rect 48688 29504 48740 29510
rect 48688 29446 48740 29452
rect 48226 29135 48282 29144
rect 48320 29164 48372 29170
rect 48320 29106 48372 29112
rect 48136 29028 48188 29034
rect 48136 28970 48188 28976
rect 48136 28688 48188 28694
rect 48188 28636 48268 28642
rect 48136 28630 48268 28636
rect 48148 28614 48268 28630
rect 48240 28558 48268 28614
rect 48596 28620 48648 28626
rect 48596 28562 48648 28568
rect 48228 28552 48280 28558
rect 48228 28494 48280 28500
rect 47860 28076 47912 28082
rect 47860 28018 47912 28024
rect 48044 28076 48096 28082
rect 48044 28018 48096 28024
rect 47872 27470 47900 28018
rect 47952 27872 48004 27878
rect 47952 27814 48004 27820
rect 47964 27713 47992 27814
rect 47950 27704 48006 27713
rect 47950 27639 48006 27648
rect 47860 27464 47912 27470
rect 47860 27406 47912 27412
rect 47964 27402 47992 27639
rect 48056 27538 48084 28018
rect 48044 27532 48096 27538
rect 48044 27474 48096 27480
rect 47952 27396 48004 27402
rect 47952 27338 48004 27344
rect 48056 27130 48084 27474
rect 48136 27464 48188 27470
rect 48136 27406 48188 27412
rect 48044 27124 48096 27130
rect 48044 27066 48096 27072
rect 48148 26994 48176 27406
rect 48608 27402 48636 28562
rect 48596 27396 48648 27402
rect 48596 27338 48648 27344
rect 48136 26988 48188 26994
rect 48136 26930 48188 26936
rect 48148 26790 48176 26930
rect 48136 26784 48188 26790
rect 48136 26726 48188 26732
rect 48148 26382 48176 26726
rect 48228 26444 48280 26450
rect 48228 26386 48280 26392
rect 48136 26376 48188 26382
rect 48136 26318 48188 26324
rect 48240 25906 48268 26386
rect 48320 26308 48372 26314
rect 48700 26296 48728 29446
rect 48780 28960 48832 28966
rect 48780 28902 48832 28908
rect 48792 28082 48820 28902
rect 48884 28694 48912 30194
rect 49160 30190 49188 30246
rect 49148 30184 49200 30190
rect 49148 30126 49200 30132
rect 49160 29850 49188 30126
rect 49148 29844 49200 29850
rect 49148 29786 49200 29792
rect 49056 29776 49108 29782
rect 49056 29718 49108 29724
rect 48872 28688 48924 28694
rect 48872 28630 48924 28636
rect 48780 28076 48832 28082
rect 48780 28018 48832 28024
rect 48884 27606 48912 28630
rect 49068 28558 49096 29718
rect 49424 29572 49476 29578
rect 49424 29514 49476 29520
rect 49148 28960 49200 28966
rect 49148 28902 49200 28908
rect 49332 28960 49384 28966
rect 49332 28902 49384 28908
rect 49160 28626 49188 28902
rect 49344 28762 49372 28902
rect 49332 28756 49384 28762
rect 49332 28698 49384 28704
rect 49148 28620 49200 28626
rect 49148 28562 49200 28568
rect 49436 28558 49464 29514
rect 49712 29510 49740 30262
rect 49700 29504 49752 29510
rect 49700 29446 49752 29452
rect 49792 29504 49844 29510
rect 49792 29446 49844 29452
rect 49516 29164 49568 29170
rect 49700 29164 49752 29170
rect 49568 29124 49648 29152
rect 49516 29106 49568 29112
rect 49620 28642 49648 29124
rect 49700 29106 49752 29112
rect 49712 28762 49740 29106
rect 49700 28756 49752 28762
rect 49700 28698 49752 28704
rect 49620 28614 49740 28642
rect 49056 28552 49108 28558
rect 49056 28494 49108 28500
rect 49424 28552 49476 28558
rect 49476 28512 49556 28540
rect 49424 28494 49476 28500
rect 49332 28416 49384 28422
rect 49332 28358 49384 28364
rect 48962 28112 49018 28121
rect 48962 28047 48964 28056
rect 49016 28047 49018 28056
rect 48964 28018 49016 28024
rect 48872 27600 48924 27606
rect 48872 27542 48924 27548
rect 48884 26926 48912 27542
rect 48964 26988 49016 26994
rect 48964 26930 49016 26936
rect 48872 26920 48924 26926
rect 48872 26862 48924 26868
rect 48872 26512 48924 26518
rect 48872 26454 48924 26460
rect 48780 26308 48832 26314
rect 48700 26268 48780 26296
rect 48320 26250 48372 26256
rect 48780 26250 48832 26256
rect 48228 25900 48280 25906
rect 48228 25842 48280 25848
rect 47860 25764 47912 25770
rect 47860 25706 47912 25712
rect 47872 24818 47900 25706
rect 48240 25498 48268 25842
rect 48228 25492 48280 25498
rect 48228 25434 48280 25440
rect 48332 25294 48360 26250
rect 48412 25900 48464 25906
rect 48412 25842 48464 25848
rect 48424 25430 48452 25842
rect 48884 25702 48912 26454
rect 48976 26382 49004 26930
rect 49056 26920 49108 26926
rect 49056 26862 49108 26868
rect 48964 26376 49016 26382
rect 48964 26318 49016 26324
rect 48688 25696 48740 25702
rect 48688 25638 48740 25644
rect 48872 25696 48924 25702
rect 48872 25638 48924 25644
rect 48412 25424 48464 25430
rect 48412 25366 48464 25372
rect 48320 25288 48372 25294
rect 48320 25230 48372 25236
rect 48228 25152 48280 25158
rect 48228 25094 48280 25100
rect 47860 24812 47912 24818
rect 47860 24754 47912 24760
rect 47768 23724 47820 23730
rect 47768 23666 47820 23672
rect 47228 23186 47440 23202
rect 47216 23180 47440 23186
rect 47268 23174 47440 23180
rect 47216 23122 47268 23128
rect 47124 23044 47176 23050
rect 47124 22986 47176 22992
rect 47136 22098 47164 22986
rect 47412 22642 47440 23174
rect 47400 22636 47452 22642
rect 47400 22578 47452 22584
rect 47124 22092 47176 22098
rect 47412 22094 47440 22578
rect 47124 22034 47176 22040
rect 47320 22066 47440 22094
rect 47032 22024 47084 22030
rect 47032 21966 47084 21972
rect 39120 21684 39172 21690
rect 39120 21626 39172 21632
rect 37648 21548 37700 21554
rect 37648 21490 37700 21496
rect 38660 21548 38712 21554
rect 38660 21490 38712 21496
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 47320 21146 47348 22066
rect 47780 21690 47808 23666
rect 48240 22098 48268 25094
rect 48332 24410 48360 25230
rect 48700 24682 48728 25638
rect 48780 24812 48832 24818
rect 48780 24754 48832 24760
rect 48688 24676 48740 24682
rect 48688 24618 48740 24624
rect 48320 24404 48372 24410
rect 48320 24346 48372 24352
rect 48792 23730 48820 24754
rect 48780 23724 48832 23730
rect 48780 23666 48832 23672
rect 48884 23186 48912 25638
rect 49068 25498 49096 26862
rect 49344 26382 49372 28358
rect 49528 27538 49556 28512
rect 49606 28248 49662 28257
rect 49712 28218 49740 28614
rect 49606 28183 49608 28192
rect 49660 28183 49662 28192
rect 49700 28212 49752 28218
rect 49608 28154 49660 28160
rect 49700 28154 49752 28160
rect 49608 28008 49660 28014
rect 49608 27950 49660 27956
rect 49620 27606 49648 27950
rect 49712 27690 49740 28154
rect 49804 27878 49832 29446
rect 49896 29306 49924 31078
rect 50172 29646 50200 39850
rect 50712 38956 50764 38962
rect 50712 38898 50764 38904
rect 50344 38752 50396 38758
rect 50344 38694 50396 38700
rect 50356 38350 50384 38694
rect 50344 38344 50396 38350
rect 50344 38286 50396 38292
rect 50436 38344 50488 38350
rect 50436 38286 50488 38292
rect 50448 37670 50476 38286
rect 50724 38282 50752 38898
rect 50816 38826 50844 41074
rect 50908 40594 50936 41414
rect 50896 40588 50948 40594
rect 50896 40530 50948 40536
rect 51000 39370 51028 41414
rect 51092 41274 51120 41754
rect 51172 41608 51224 41614
rect 51172 41550 51224 41556
rect 51080 41268 51132 41274
rect 51080 41210 51132 41216
rect 51184 40934 51212 41550
rect 51172 40928 51224 40934
rect 51172 40870 51224 40876
rect 51172 40588 51224 40594
rect 51172 40530 51224 40536
rect 51184 40390 51212 40530
rect 51460 40474 51488 43182
rect 51724 42560 51776 42566
rect 51724 42502 51776 42508
rect 51736 42090 51764 42502
rect 51724 42084 51776 42090
rect 51724 42026 51776 42032
rect 51540 41676 51592 41682
rect 51540 41618 51592 41624
rect 51552 40662 51580 41618
rect 51724 41472 51776 41478
rect 51724 41414 51776 41420
rect 51736 41206 51764 41414
rect 51724 41200 51776 41206
rect 51724 41142 51776 41148
rect 51828 41138 51856 43726
rect 52012 42702 52040 44882
rect 52104 44470 52132 45766
rect 53012 44940 53064 44946
rect 53012 44882 53064 44888
rect 52644 44736 52696 44742
rect 52644 44678 52696 44684
rect 52092 44464 52144 44470
rect 52092 44406 52144 44412
rect 52104 43654 52132 44406
rect 52276 44260 52328 44266
rect 52276 44202 52328 44208
rect 52092 43648 52144 43654
rect 52092 43590 52144 43596
rect 52104 43450 52132 43590
rect 52092 43444 52144 43450
rect 52092 43386 52144 43392
rect 52000 42696 52052 42702
rect 52000 42638 52052 42644
rect 52012 42537 52040 42638
rect 51998 42528 52054 42537
rect 51998 42463 52054 42472
rect 52092 42152 52144 42158
rect 52092 42094 52144 42100
rect 52104 41750 52132 42094
rect 52184 42016 52236 42022
rect 52184 41958 52236 41964
rect 51908 41744 51960 41750
rect 51908 41686 51960 41692
rect 52092 41744 52144 41750
rect 52092 41686 52144 41692
rect 51920 41206 51948 41686
rect 52000 41472 52052 41478
rect 52000 41414 52052 41420
rect 51908 41200 51960 41206
rect 51908 41142 51960 41148
rect 52012 41138 52040 41414
rect 51632 41132 51684 41138
rect 51632 41074 51684 41080
rect 51816 41132 51868 41138
rect 51816 41074 51868 41080
rect 52000 41132 52052 41138
rect 52000 41074 52052 41080
rect 51540 40656 51592 40662
rect 51540 40598 51592 40604
rect 51264 40452 51316 40458
rect 51460 40446 51580 40474
rect 51264 40394 51316 40400
rect 51172 40384 51224 40390
rect 51172 40326 51224 40332
rect 50988 39364 51040 39370
rect 50988 39306 51040 39312
rect 51080 38956 51132 38962
rect 51080 38898 51132 38904
rect 50804 38820 50856 38826
rect 50804 38762 50856 38768
rect 51092 38554 51120 38898
rect 51172 38888 51224 38894
rect 51172 38830 51224 38836
rect 51080 38548 51132 38554
rect 51080 38490 51132 38496
rect 51184 38486 51212 38830
rect 51172 38480 51224 38486
rect 50802 38448 50858 38457
rect 51172 38422 51224 38428
rect 50802 38383 50858 38392
rect 50816 38350 50844 38383
rect 50804 38344 50856 38350
rect 50804 38286 50856 38292
rect 50712 38276 50764 38282
rect 50712 38218 50764 38224
rect 50896 38276 50948 38282
rect 50896 38218 50948 38224
rect 50436 37664 50488 37670
rect 50436 37606 50488 37612
rect 50252 37324 50304 37330
rect 50252 37266 50304 37272
rect 50264 35698 50292 37266
rect 50344 37188 50396 37194
rect 50344 37130 50396 37136
rect 50356 36854 50384 37130
rect 50724 36922 50752 38218
rect 50804 37800 50856 37806
rect 50804 37742 50856 37748
rect 50816 37262 50844 37742
rect 50908 37670 50936 38218
rect 50896 37664 50948 37670
rect 50896 37606 50948 37612
rect 50804 37256 50856 37262
rect 50804 37198 50856 37204
rect 50988 37256 51040 37262
rect 50988 37198 51040 37204
rect 50712 36916 50764 36922
rect 50712 36858 50764 36864
rect 50344 36848 50396 36854
rect 50344 36790 50396 36796
rect 50344 36576 50396 36582
rect 50344 36518 50396 36524
rect 50712 36576 50764 36582
rect 50712 36518 50764 36524
rect 50356 36174 50384 36518
rect 50724 36310 50752 36518
rect 50712 36304 50764 36310
rect 50712 36246 50764 36252
rect 50344 36168 50396 36174
rect 50344 36110 50396 36116
rect 50620 36168 50672 36174
rect 50620 36110 50672 36116
rect 50632 35766 50660 36110
rect 50620 35760 50672 35766
rect 50620 35702 50672 35708
rect 50724 35698 50752 36246
rect 51000 36242 51028 37198
rect 50988 36236 51040 36242
rect 50988 36178 51040 36184
rect 51276 36174 51304 40394
rect 51448 40384 51500 40390
rect 51448 40326 51500 40332
rect 50896 36168 50948 36174
rect 50896 36110 50948 36116
rect 51264 36168 51316 36174
rect 51264 36110 51316 36116
rect 50804 36032 50856 36038
rect 50804 35974 50856 35980
rect 50252 35692 50304 35698
rect 50252 35634 50304 35640
rect 50712 35692 50764 35698
rect 50712 35634 50764 35640
rect 50620 35624 50672 35630
rect 50620 35566 50672 35572
rect 50632 34134 50660 35566
rect 50724 34932 50752 35634
rect 50816 35086 50844 35974
rect 50908 35562 50936 36110
rect 50988 35828 51040 35834
rect 50988 35770 51040 35776
rect 50896 35556 50948 35562
rect 50896 35498 50948 35504
rect 50804 35080 50856 35086
rect 50804 35022 50856 35028
rect 50724 34904 50844 34932
rect 50816 34610 50844 34904
rect 51000 34746 51028 35770
rect 51356 34944 51408 34950
rect 51356 34886 51408 34892
rect 50988 34740 51040 34746
rect 50988 34682 51040 34688
rect 50804 34604 50856 34610
rect 50804 34546 50856 34552
rect 50620 34128 50672 34134
rect 50620 34070 50672 34076
rect 50252 33856 50304 33862
rect 50252 33798 50304 33804
rect 50264 33522 50292 33798
rect 50252 33516 50304 33522
rect 50252 33458 50304 33464
rect 50816 33114 50844 34546
rect 50988 33992 51040 33998
rect 50988 33934 51040 33940
rect 51000 33454 51028 33934
rect 51368 33930 51396 34886
rect 51460 34610 51488 40326
rect 51448 34604 51500 34610
rect 51448 34546 51500 34552
rect 51552 34542 51580 40446
rect 51644 39370 51672 41074
rect 51724 39840 51776 39846
rect 51724 39782 51776 39788
rect 51736 39506 51764 39782
rect 51724 39500 51776 39506
rect 51724 39442 51776 39448
rect 51828 39438 51856 41074
rect 52000 40928 52052 40934
rect 52000 40870 52052 40876
rect 52012 40526 52040 40870
rect 52104 40526 52132 41686
rect 52196 41614 52224 41958
rect 52184 41608 52236 41614
rect 52184 41550 52236 41556
rect 52288 41546 52316 44202
rect 52656 44198 52684 44678
rect 53024 44402 53052 44882
rect 52828 44396 52880 44402
rect 52828 44338 52880 44344
rect 53012 44396 53064 44402
rect 53012 44338 53064 44344
rect 54576 44396 54628 44402
rect 54576 44338 54628 44344
rect 55772 44396 55824 44402
rect 55772 44338 55824 44344
rect 52644 44192 52696 44198
rect 52644 44134 52696 44140
rect 52656 43110 52684 44134
rect 52840 43178 52868 44338
rect 54588 43994 54616 44338
rect 54576 43988 54628 43994
rect 54576 43930 54628 43936
rect 53932 43920 53984 43926
rect 53932 43862 53984 43868
rect 53656 43784 53708 43790
rect 53656 43726 53708 43732
rect 53288 43648 53340 43654
rect 53288 43590 53340 43596
rect 52828 43172 52880 43178
rect 52828 43114 52880 43120
rect 52644 43104 52696 43110
rect 52644 43046 52696 43052
rect 52656 42362 52684 43046
rect 52460 42356 52512 42362
rect 52460 42298 52512 42304
rect 52644 42356 52696 42362
rect 52644 42298 52696 42304
rect 52276 41540 52328 41546
rect 52276 41482 52328 41488
rect 52000 40520 52052 40526
rect 52000 40462 52052 40468
rect 52092 40520 52144 40526
rect 52092 40462 52144 40468
rect 52104 40050 52132 40462
rect 52288 40458 52316 41482
rect 52368 41132 52420 41138
rect 52368 41074 52420 41080
rect 52380 40526 52408 41074
rect 52368 40520 52420 40526
rect 52368 40462 52420 40468
rect 52276 40452 52328 40458
rect 52276 40394 52328 40400
rect 52092 40044 52144 40050
rect 52092 39986 52144 39992
rect 52104 39574 52132 39986
rect 52092 39568 52144 39574
rect 52092 39510 52144 39516
rect 51816 39432 51868 39438
rect 51816 39374 51868 39380
rect 51632 39364 51684 39370
rect 51632 39306 51684 39312
rect 51644 39030 51672 39306
rect 51724 39296 51776 39302
rect 51724 39238 51776 39244
rect 51736 39030 51764 39238
rect 51632 39024 51684 39030
rect 51632 38966 51684 38972
rect 51724 39024 51776 39030
rect 51724 38966 51776 38972
rect 51828 38826 51856 39374
rect 51908 39296 51960 39302
rect 51908 39238 51960 39244
rect 51920 38944 51948 39238
rect 52000 38956 52052 38962
rect 51920 38916 52000 38944
rect 51816 38820 51868 38826
rect 51816 38762 51868 38768
rect 51920 38554 51948 38916
rect 52000 38898 52052 38904
rect 52288 38826 52316 40394
rect 52000 38820 52052 38826
rect 52000 38762 52052 38768
rect 52276 38820 52328 38826
rect 52276 38762 52328 38768
rect 51908 38548 51960 38554
rect 51908 38490 51960 38496
rect 51920 38010 51948 38490
rect 52012 38214 52040 38762
rect 52380 38282 52408 40462
rect 52368 38276 52420 38282
rect 52368 38218 52420 38224
rect 52000 38208 52052 38214
rect 52000 38150 52052 38156
rect 51908 38004 51960 38010
rect 51908 37946 51960 37952
rect 52368 38004 52420 38010
rect 52368 37946 52420 37952
rect 52000 37392 52052 37398
rect 52000 37334 52052 37340
rect 52012 37126 52040 37334
rect 52000 37120 52052 37126
rect 52000 37062 52052 37068
rect 52012 36854 52040 37062
rect 52380 36922 52408 37946
rect 52472 37618 52500 42298
rect 52656 41682 52684 42298
rect 52644 41676 52696 41682
rect 52644 41618 52696 41624
rect 52472 37590 52592 37618
rect 52460 37460 52512 37466
rect 52460 37402 52512 37408
rect 52472 37194 52500 37402
rect 52460 37188 52512 37194
rect 52460 37130 52512 37136
rect 52368 36916 52420 36922
rect 52368 36858 52420 36864
rect 52000 36848 52052 36854
rect 51920 36796 52000 36802
rect 51920 36790 52052 36796
rect 51920 36774 52040 36790
rect 52092 36780 52144 36786
rect 51632 36032 51684 36038
rect 51632 35974 51684 35980
rect 51540 34536 51592 34542
rect 51540 34478 51592 34484
rect 51644 34134 51672 35974
rect 51920 35494 51948 36774
rect 52092 36722 52144 36728
rect 52276 36780 52328 36786
rect 52276 36722 52328 36728
rect 52104 36038 52132 36722
rect 52092 36032 52144 36038
rect 52092 35974 52144 35980
rect 51908 35488 51960 35494
rect 51908 35430 51960 35436
rect 51724 34604 51776 34610
rect 51724 34546 51776 34552
rect 51632 34128 51684 34134
rect 51632 34070 51684 34076
rect 51356 33924 51408 33930
rect 51356 33866 51408 33872
rect 51644 33862 51672 34070
rect 51632 33856 51684 33862
rect 51632 33798 51684 33804
rect 51356 33516 51408 33522
rect 51356 33458 51408 33464
rect 50988 33448 51040 33454
rect 50988 33390 51040 33396
rect 51080 33448 51132 33454
rect 51080 33390 51132 33396
rect 50804 33108 50856 33114
rect 50804 33050 50856 33056
rect 50712 32836 50764 32842
rect 50712 32778 50764 32784
rect 50724 32434 50752 32778
rect 50816 32570 50844 33050
rect 51092 32978 51120 33390
rect 51080 32972 51132 32978
rect 51080 32914 51132 32920
rect 51368 32570 51396 33458
rect 51632 32836 51684 32842
rect 51632 32778 51684 32784
rect 50804 32564 50856 32570
rect 50804 32506 50856 32512
rect 51356 32564 51408 32570
rect 51356 32506 51408 32512
rect 50712 32428 50764 32434
rect 50712 32370 50764 32376
rect 50816 31754 50844 32506
rect 51644 32434 51672 32778
rect 50896 32428 50948 32434
rect 50896 32370 50948 32376
rect 51080 32428 51132 32434
rect 51080 32370 51132 32376
rect 51632 32428 51684 32434
rect 51632 32370 51684 32376
rect 50908 31890 50936 32370
rect 50988 32360 51040 32366
rect 50988 32302 51040 32308
rect 50896 31884 50948 31890
rect 50896 31826 50948 31832
rect 51000 31822 51028 32302
rect 50988 31816 51040 31822
rect 50988 31758 51040 31764
rect 50804 31748 50856 31754
rect 50804 31690 50856 31696
rect 50816 31346 50844 31690
rect 50988 31476 51040 31482
rect 51092 31464 51120 32370
rect 51448 31816 51500 31822
rect 51448 31758 51500 31764
rect 51632 31816 51684 31822
rect 51632 31758 51684 31764
rect 51040 31436 51120 31464
rect 50988 31418 51040 31424
rect 50804 31340 50856 31346
rect 50804 31282 50856 31288
rect 50344 31204 50396 31210
rect 50344 31146 50396 31152
rect 50356 30802 50384 31146
rect 51356 31136 51408 31142
rect 51356 31078 51408 31084
rect 50988 30864 51040 30870
rect 50988 30806 51040 30812
rect 50344 30796 50396 30802
rect 50344 30738 50396 30744
rect 50804 30796 50856 30802
rect 50804 30738 50856 30744
rect 50620 30660 50672 30666
rect 50620 30602 50672 30608
rect 50632 30326 50660 30602
rect 50436 30320 50488 30326
rect 50620 30320 50672 30326
rect 50488 30280 50620 30308
rect 50436 30262 50488 30268
rect 50620 30262 50672 30268
rect 50252 30048 50304 30054
rect 50252 29990 50304 29996
rect 50160 29640 50212 29646
rect 50160 29582 50212 29588
rect 49884 29300 49936 29306
rect 49884 29242 49936 29248
rect 49896 29170 49924 29242
rect 50172 29238 50200 29582
rect 50160 29232 50212 29238
rect 50160 29174 50212 29180
rect 49884 29164 49936 29170
rect 49884 29106 49936 29112
rect 50264 28014 50292 29990
rect 50342 29200 50398 29209
rect 50632 29170 50660 30262
rect 50816 30258 50844 30738
rect 50804 30252 50856 30258
rect 50804 30194 50856 30200
rect 50342 29135 50398 29144
rect 50620 29164 50672 29170
rect 50356 28558 50384 29135
rect 50620 29106 50672 29112
rect 50804 28960 50856 28966
rect 50804 28902 50856 28908
rect 50816 28694 50844 28902
rect 50436 28688 50488 28694
rect 50804 28688 50856 28694
rect 50488 28636 50660 28642
rect 50436 28630 50660 28636
rect 50804 28630 50856 28636
rect 50448 28614 50660 28630
rect 50632 28558 50660 28614
rect 50344 28552 50396 28558
rect 50344 28494 50396 28500
rect 50528 28552 50580 28558
rect 50528 28494 50580 28500
rect 50620 28552 50672 28558
rect 50620 28494 50672 28500
rect 50540 28218 50568 28494
rect 50528 28212 50580 28218
rect 50528 28154 50580 28160
rect 50344 28144 50396 28150
rect 50344 28086 50396 28092
rect 50252 28008 50304 28014
rect 50252 27950 50304 27956
rect 49792 27872 49844 27878
rect 49792 27814 49844 27820
rect 49712 27662 49832 27690
rect 49608 27600 49660 27606
rect 49608 27542 49660 27548
rect 49516 27532 49568 27538
rect 49516 27474 49568 27480
rect 49332 26376 49384 26382
rect 49332 26318 49384 26324
rect 49528 26042 49556 27474
rect 49608 27464 49660 27470
rect 49608 27406 49660 27412
rect 49620 26790 49648 27406
rect 49804 27334 49832 27662
rect 49884 27668 49936 27674
rect 49884 27610 49936 27616
rect 49792 27328 49844 27334
rect 49792 27270 49844 27276
rect 49608 26784 49660 26790
rect 49608 26726 49660 26732
rect 49620 26382 49648 26726
rect 49700 26444 49752 26450
rect 49700 26386 49752 26392
rect 49608 26376 49660 26382
rect 49608 26318 49660 26324
rect 49516 26036 49568 26042
rect 49516 25978 49568 25984
rect 49056 25492 49108 25498
rect 49056 25434 49108 25440
rect 49620 25294 49648 26318
rect 49712 25344 49740 26386
rect 49804 25906 49832 27270
rect 49896 25906 49924 27610
rect 50356 26994 50384 28086
rect 50620 28076 50672 28082
rect 50620 28018 50672 28024
rect 50436 28008 50488 28014
rect 50436 27950 50488 27956
rect 50448 27674 50476 27950
rect 50528 27872 50580 27878
rect 50528 27814 50580 27820
rect 50436 27668 50488 27674
rect 50436 27610 50488 27616
rect 50436 27464 50488 27470
rect 50436 27406 50488 27412
rect 50068 26988 50120 26994
rect 50068 26930 50120 26936
rect 50160 26988 50212 26994
rect 50160 26930 50212 26936
rect 50344 26988 50396 26994
rect 50344 26930 50396 26936
rect 49792 25900 49844 25906
rect 49792 25842 49844 25848
rect 49884 25900 49936 25906
rect 49884 25842 49936 25848
rect 50080 25362 50108 26930
rect 50172 25974 50200 26930
rect 50160 25968 50212 25974
rect 50160 25910 50212 25916
rect 49884 25356 49936 25362
rect 49712 25316 49832 25344
rect 49608 25288 49660 25294
rect 49608 25230 49660 25236
rect 49620 24274 49648 25230
rect 49700 25220 49752 25226
rect 49700 25162 49752 25168
rect 49608 24268 49660 24274
rect 49608 24210 49660 24216
rect 49712 24206 49740 25162
rect 49700 24200 49752 24206
rect 49700 24142 49752 24148
rect 49056 24132 49108 24138
rect 49056 24074 49108 24080
rect 49068 23866 49096 24074
rect 49056 23860 49108 23866
rect 49056 23802 49108 23808
rect 49148 23724 49200 23730
rect 49148 23666 49200 23672
rect 49160 23526 49188 23666
rect 49148 23520 49200 23526
rect 49148 23462 49200 23468
rect 48872 23180 48924 23186
rect 48872 23122 48924 23128
rect 48320 22568 48372 22574
rect 48320 22510 48372 22516
rect 48332 22234 48360 22510
rect 48320 22228 48372 22234
rect 48320 22170 48372 22176
rect 49160 22098 49188 23462
rect 49712 22778 49740 24142
rect 49804 23798 49832 25316
rect 49884 25298 49936 25304
rect 50068 25356 50120 25362
rect 50068 25298 50120 25304
rect 49896 24070 49924 25298
rect 50172 25294 50200 25910
rect 50160 25288 50212 25294
rect 50160 25230 50212 25236
rect 50252 24608 50304 24614
rect 50252 24550 50304 24556
rect 49884 24064 49936 24070
rect 49884 24006 49936 24012
rect 49792 23792 49844 23798
rect 49792 23734 49844 23740
rect 49804 23118 49832 23734
rect 49884 23656 49936 23662
rect 49884 23598 49936 23604
rect 49896 23254 49924 23598
rect 49884 23248 49936 23254
rect 49884 23190 49936 23196
rect 50264 23118 50292 24550
rect 50356 24410 50384 26930
rect 50448 26364 50476 27406
rect 50540 26994 50568 27814
rect 50632 27470 50660 28018
rect 50620 27464 50672 27470
rect 50620 27406 50672 27412
rect 50528 26988 50580 26994
rect 50528 26930 50580 26936
rect 50632 26586 50660 27406
rect 50620 26580 50672 26586
rect 50620 26522 50672 26528
rect 50528 26376 50580 26382
rect 50448 26336 50528 26364
rect 50528 26318 50580 26324
rect 50540 26246 50568 26318
rect 50528 26240 50580 26246
rect 50528 26182 50580 26188
rect 50816 25974 50844 28630
rect 50896 27328 50948 27334
rect 50896 27270 50948 27276
rect 50908 26926 50936 27270
rect 50896 26920 50948 26926
rect 50896 26862 50948 26868
rect 51000 26246 51028 30806
rect 51172 30728 51224 30734
rect 51172 30670 51224 30676
rect 51184 30394 51212 30670
rect 51172 30388 51224 30394
rect 51172 30330 51224 30336
rect 51368 29170 51396 31078
rect 51460 30802 51488 31758
rect 51540 31340 51592 31346
rect 51540 31282 51592 31288
rect 51552 30938 51580 31282
rect 51540 30932 51592 30938
rect 51540 30874 51592 30880
rect 51448 30796 51500 30802
rect 51448 30738 51500 30744
rect 51644 30734 51672 31758
rect 51632 30728 51684 30734
rect 51632 30670 51684 30676
rect 51736 29170 51764 34546
rect 51920 32552 51948 35430
rect 52104 34202 52132 35974
rect 52288 35834 52316 36722
rect 52276 35828 52328 35834
rect 52276 35770 52328 35776
rect 52564 35290 52592 37590
rect 52552 35284 52604 35290
rect 52552 35226 52604 35232
rect 52368 34672 52420 34678
rect 52368 34614 52420 34620
rect 52092 34196 52144 34202
rect 52092 34138 52144 34144
rect 52092 33992 52144 33998
rect 52092 33934 52144 33940
rect 52000 33856 52052 33862
rect 52000 33798 52052 33804
rect 52012 33590 52040 33798
rect 52000 33584 52052 33590
rect 52000 33526 52052 33532
rect 52000 32564 52052 32570
rect 51920 32524 52000 32552
rect 52000 32506 52052 32512
rect 52012 32434 52040 32506
rect 51908 32428 51960 32434
rect 51908 32370 51960 32376
rect 52000 32428 52052 32434
rect 52000 32370 52052 32376
rect 51920 31958 51948 32370
rect 51908 31952 51960 31958
rect 51908 31894 51960 31900
rect 51920 31414 51948 31894
rect 51908 31408 51960 31414
rect 51908 31350 51960 31356
rect 52000 30660 52052 30666
rect 52000 30602 52052 30608
rect 52012 30258 52040 30602
rect 52000 30252 52052 30258
rect 52000 30194 52052 30200
rect 51908 30048 51960 30054
rect 51908 29990 51960 29996
rect 51920 29714 51948 29990
rect 51908 29708 51960 29714
rect 51908 29650 51960 29656
rect 52104 29646 52132 33934
rect 52380 33522 52408 34614
rect 52460 34468 52512 34474
rect 52460 34410 52512 34416
rect 52472 33590 52500 34410
rect 52460 33584 52512 33590
rect 52460 33526 52512 33532
rect 52368 33516 52420 33522
rect 52368 33458 52420 33464
rect 52380 33114 52408 33458
rect 52368 33108 52420 33114
rect 52368 33050 52420 33056
rect 52276 32972 52328 32978
rect 52276 32914 52328 32920
rect 52184 32428 52236 32434
rect 52184 32370 52236 32376
rect 52196 32026 52224 32370
rect 52288 32298 52316 32914
rect 52564 32910 52592 35226
rect 52656 34950 52684 41618
rect 52840 41614 52868 43114
rect 53300 42702 53328 43590
rect 53472 43104 53524 43110
rect 53472 43046 53524 43052
rect 53380 42764 53432 42770
rect 53380 42706 53432 42712
rect 53104 42696 53156 42702
rect 53104 42638 53156 42644
rect 53288 42696 53340 42702
rect 53288 42638 53340 42644
rect 53116 42362 53144 42638
rect 53104 42356 53156 42362
rect 53104 42298 53156 42304
rect 53012 42220 53064 42226
rect 53012 42162 53064 42168
rect 52828 41608 52880 41614
rect 52828 41550 52880 41556
rect 52840 40458 52868 41550
rect 53024 40746 53052 42162
rect 53392 42158 53420 42706
rect 53484 42702 53512 43046
rect 53668 42906 53696 43726
rect 53944 43450 53972 43862
rect 55496 43852 55548 43858
rect 55496 43794 55548 43800
rect 55312 43784 55364 43790
rect 55312 43726 55364 43732
rect 55036 43716 55088 43722
rect 55036 43658 55088 43664
rect 54484 43648 54536 43654
rect 54484 43590 54536 43596
rect 53932 43444 53984 43450
rect 53932 43386 53984 43392
rect 54300 43444 54352 43450
rect 54300 43386 54352 43392
rect 53656 42900 53708 42906
rect 53656 42842 53708 42848
rect 54312 42770 54340 43386
rect 54300 42764 54352 42770
rect 54300 42706 54352 42712
rect 53472 42696 53524 42702
rect 53472 42638 53524 42644
rect 53656 42696 53708 42702
rect 53656 42638 53708 42644
rect 53668 42294 53696 42638
rect 53748 42628 53800 42634
rect 53748 42570 53800 42576
rect 53656 42288 53708 42294
rect 53656 42230 53708 42236
rect 53760 42226 53788 42570
rect 53932 42560 53984 42566
rect 53932 42502 53984 42508
rect 53748 42220 53800 42226
rect 53748 42162 53800 42168
rect 53944 42158 53972 42502
rect 54312 42226 54340 42706
rect 54392 42696 54444 42702
rect 54392 42638 54444 42644
rect 54116 42220 54168 42226
rect 54116 42162 54168 42168
rect 54300 42220 54352 42226
rect 54300 42162 54352 42168
rect 53196 42152 53248 42158
rect 53196 42094 53248 42100
rect 53380 42152 53432 42158
rect 53380 42094 53432 42100
rect 53932 42152 53984 42158
rect 53932 42094 53984 42100
rect 53104 42016 53156 42022
rect 53104 41958 53156 41964
rect 53116 41682 53144 41958
rect 53104 41676 53156 41682
rect 53104 41618 53156 41624
rect 53104 40928 53156 40934
rect 53104 40870 53156 40876
rect 52932 40718 53052 40746
rect 52828 40452 52880 40458
rect 52828 40394 52880 40400
rect 52840 38962 52868 40394
rect 52932 39982 52960 40718
rect 53116 40390 53144 40870
rect 53104 40384 53156 40390
rect 53104 40326 53156 40332
rect 52920 39976 52972 39982
rect 52920 39918 52972 39924
rect 52828 38956 52880 38962
rect 52828 38898 52880 38904
rect 52736 38752 52788 38758
rect 52736 38694 52788 38700
rect 52748 36174 52776 38694
rect 52840 38457 52868 38898
rect 52932 38554 52960 39918
rect 53208 39914 53236 42094
rect 53564 41676 53616 41682
rect 53564 41618 53616 41624
rect 53380 40520 53432 40526
rect 53380 40462 53432 40468
rect 53392 40118 53420 40462
rect 53576 40118 53604 41618
rect 53944 41614 53972 42094
rect 54024 42016 54076 42022
rect 54024 41958 54076 41964
rect 54036 41682 54064 41958
rect 54024 41676 54076 41682
rect 54024 41618 54076 41624
rect 53932 41608 53984 41614
rect 53932 41550 53984 41556
rect 53840 41472 53892 41478
rect 53840 41414 53892 41420
rect 53852 41138 53880 41414
rect 53840 41132 53892 41138
rect 53840 41074 53892 41080
rect 53944 40934 53972 41550
rect 54024 41132 54076 41138
rect 54024 41074 54076 41080
rect 53932 40928 53984 40934
rect 53852 40888 53932 40916
rect 53852 40594 53880 40888
rect 53932 40870 53984 40876
rect 54036 40610 54064 41074
rect 54128 40730 54156 42162
rect 54312 41478 54340 42162
rect 54404 42022 54432 42638
rect 54496 42566 54524 43590
rect 54944 43308 54996 43314
rect 54944 43250 54996 43256
rect 54956 42906 54984 43250
rect 54944 42900 54996 42906
rect 54944 42842 54996 42848
rect 54760 42764 54812 42770
rect 54760 42706 54812 42712
rect 54484 42560 54536 42566
rect 54484 42502 54536 42508
rect 54772 42362 54800 42706
rect 54760 42356 54812 42362
rect 54760 42298 54812 42304
rect 55048 42294 55076 43658
rect 55324 43246 55352 43726
rect 55312 43240 55364 43246
rect 55312 43182 55364 43188
rect 55220 43172 55272 43178
rect 55220 43114 55272 43120
rect 55128 43104 55180 43110
rect 55128 43046 55180 43052
rect 55140 42702 55168 43046
rect 55232 42838 55260 43114
rect 55220 42832 55272 42838
rect 55220 42774 55272 42780
rect 55128 42696 55180 42702
rect 55128 42638 55180 42644
rect 55140 42362 55168 42638
rect 55128 42356 55180 42362
rect 55128 42298 55180 42304
rect 55036 42288 55088 42294
rect 55036 42230 55088 42236
rect 54576 42220 54628 42226
rect 54576 42162 54628 42168
rect 54392 42016 54444 42022
rect 54392 41958 54444 41964
rect 54392 41540 54444 41546
rect 54392 41482 54444 41488
rect 54300 41472 54352 41478
rect 54300 41414 54352 41420
rect 54404 41206 54432 41482
rect 54484 41472 54536 41478
rect 54484 41414 54536 41420
rect 54392 41200 54444 41206
rect 54392 41142 54444 41148
rect 54496 41070 54524 41414
rect 54484 41064 54536 41070
rect 54484 41006 54536 41012
rect 54588 41002 54616 42162
rect 55048 42158 55076 42230
rect 55036 42152 55088 42158
rect 55036 42094 55088 42100
rect 55048 41478 55076 42094
rect 55036 41472 55088 41478
rect 55036 41414 55088 41420
rect 54760 41200 54812 41206
rect 54760 41142 54812 41148
rect 54668 41064 54720 41070
rect 54668 41006 54720 41012
rect 54576 40996 54628 41002
rect 54576 40938 54628 40944
rect 54116 40724 54168 40730
rect 54116 40666 54168 40672
rect 53656 40588 53708 40594
rect 53656 40530 53708 40536
rect 53840 40588 53892 40594
rect 54036 40582 54248 40610
rect 53840 40530 53892 40536
rect 53380 40112 53432 40118
rect 53380 40054 53432 40060
rect 53564 40112 53616 40118
rect 53564 40054 53616 40060
rect 53196 39908 53248 39914
rect 53196 39850 53248 39856
rect 53392 39846 53420 40054
rect 53668 40050 53696 40530
rect 53932 40520 53984 40526
rect 53932 40462 53984 40468
rect 54024 40520 54076 40526
rect 54024 40462 54076 40468
rect 53944 40186 53972 40462
rect 54036 40202 54064 40462
rect 54036 40186 54156 40202
rect 53932 40180 53984 40186
rect 53932 40122 53984 40128
rect 54036 40180 54168 40186
rect 54036 40174 54116 40180
rect 54036 40066 54064 40174
rect 54116 40122 54168 40128
rect 53656 40044 53708 40050
rect 53656 39986 53708 39992
rect 53944 40038 54064 40066
rect 54116 40044 54168 40050
rect 53668 39930 53696 39986
rect 53564 39908 53616 39914
rect 53668 39902 53788 39930
rect 53564 39850 53616 39856
rect 53380 39840 53432 39846
rect 53380 39782 53432 39788
rect 53392 39506 53420 39782
rect 53380 39500 53432 39506
rect 53380 39442 53432 39448
rect 53012 38752 53064 38758
rect 53012 38694 53064 38700
rect 52920 38548 52972 38554
rect 52920 38490 52972 38496
rect 52826 38448 52882 38457
rect 53024 38418 53052 38694
rect 52826 38383 52882 38392
rect 53012 38412 53064 38418
rect 53012 38354 53064 38360
rect 53196 38344 53248 38350
rect 53196 38286 53248 38292
rect 53208 37874 53236 38286
rect 53196 37868 53248 37874
rect 53196 37810 53248 37816
rect 52920 37392 52972 37398
rect 52920 37334 52972 37340
rect 52932 36922 52960 37334
rect 53288 37324 53340 37330
rect 53288 37266 53340 37272
rect 53196 37120 53248 37126
rect 53196 37062 53248 37068
rect 52920 36916 52972 36922
rect 52920 36858 52972 36864
rect 52828 36576 52880 36582
rect 52828 36518 52880 36524
rect 52840 36242 52868 36518
rect 52828 36236 52880 36242
rect 52828 36178 52880 36184
rect 52736 36168 52788 36174
rect 52932 36122 52960 36858
rect 53208 36786 53236 37062
rect 53196 36780 53248 36786
rect 53196 36722 53248 36728
rect 53300 36174 53328 37266
rect 52736 36110 52788 36116
rect 52748 35698 52776 36110
rect 52840 36094 52960 36122
rect 53288 36168 53340 36174
rect 53288 36110 53340 36116
rect 52736 35692 52788 35698
rect 52736 35634 52788 35640
rect 52644 34944 52696 34950
rect 52644 34886 52696 34892
rect 52552 32904 52604 32910
rect 52552 32846 52604 32852
rect 52564 32450 52592 32846
rect 52736 32768 52788 32774
rect 52736 32710 52788 32716
rect 52748 32570 52776 32710
rect 52736 32564 52788 32570
rect 52736 32506 52788 32512
rect 52564 32434 52684 32450
rect 52564 32428 52696 32434
rect 52564 32422 52644 32428
rect 52644 32370 52696 32376
rect 52552 32360 52604 32366
rect 52552 32302 52604 32308
rect 52276 32292 52328 32298
rect 52276 32234 52328 32240
rect 52184 32020 52236 32026
rect 52184 31962 52236 31968
rect 52288 31142 52316 32234
rect 52368 32224 52420 32230
rect 52368 32166 52420 32172
rect 52380 31754 52408 32166
rect 52564 31822 52592 32302
rect 52644 32224 52696 32230
rect 52644 32166 52696 32172
rect 52552 31816 52604 31822
rect 52552 31758 52604 31764
rect 52368 31748 52420 31754
rect 52368 31690 52420 31696
rect 52656 31482 52684 32166
rect 52644 31476 52696 31482
rect 52644 31418 52696 31424
rect 52276 31136 52328 31142
rect 52276 31078 52328 31084
rect 52748 30802 52776 32506
rect 52460 30796 52512 30802
rect 52460 30738 52512 30744
rect 52736 30796 52788 30802
rect 52736 30738 52788 30744
rect 52184 30660 52236 30666
rect 52184 30602 52236 30608
rect 52196 30394 52224 30602
rect 52368 30592 52420 30598
rect 52368 30534 52420 30540
rect 52184 30388 52236 30394
rect 52184 30330 52236 30336
rect 52380 30258 52408 30534
rect 52184 30252 52236 30258
rect 52184 30194 52236 30200
rect 52368 30252 52420 30258
rect 52368 30194 52420 30200
rect 52196 30138 52224 30194
rect 52472 30138 52500 30738
rect 52552 30728 52604 30734
rect 52552 30670 52604 30676
rect 52196 30110 52500 30138
rect 52564 30122 52592 30670
rect 52840 30666 52868 36094
rect 53196 35080 53248 35086
rect 53196 35022 53248 35028
rect 52920 34604 52972 34610
rect 52920 34546 52972 34552
rect 52932 34474 52960 34546
rect 52920 34468 52972 34474
rect 52920 34410 52972 34416
rect 53012 33856 53064 33862
rect 53012 33798 53064 33804
rect 52920 32904 52972 32910
rect 52920 32846 52972 32852
rect 52932 32570 52960 32846
rect 52920 32564 52972 32570
rect 52920 32506 52972 32512
rect 52828 30660 52880 30666
rect 52828 30602 52880 30608
rect 52092 29640 52144 29646
rect 52092 29582 52144 29588
rect 51356 29164 51408 29170
rect 51356 29106 51408 29112
rect 51724 29164 51776 29170
rect 51724 29106 51776 29112
rect 51540 28960 51592 28966
rect 51540 28902 51592 28908
rect 51552 28558 51580 28902
rect 52472 28762 52500 30110
rect 52552 30116 52604 30122
rect 52552 30058 52604 30064
rect 52840 29646 52868 30602
rect 52828 29640 52880 29646
rect 52880 29588 52960 29594
rect 52828 29582 52960 29588
rect 52840 29566 52960 29582
rect 52828 29504 52880 29510
rect 52828 29446 52880 29452
rect 52840 29170 52868 29446
rect 52828 29164 52880 29170
rect 52828 29106 52880 29112
rect 52460 28756 52512 28762
rect 52460 28698 52512 28704
rect 51540 28552 51592 28558
rect 51540 28494 51592 28500
rect 52276 28552 52328 28558
rect 52276 28494 52328 28500
rect 51080 28416 51132 28422
rect 51080 28358 51132 28364
rect 51092 28121 51120 28358
rect 51998 28248 52054 28257
rect 51998 28183 52000 28192
rect 52052 28183 52054 28192
rect 52000 28154 52052 28160
rect 52288 28150 52316 28494
rect 52840 28150 52868 29106
rect 52276 28144 52328 28150
rect 51078 28112 51134 28121
rect 52276 28086 52328 28092
rect 52828 28144 52880 28150
rect 52828 28086 52880 28092
rect 51078 28047 51134 28056
rect 51356 28076 51408 28082
rect 51356 28018 51408 28024
rect 51540 28076 51592 28082
rect 51540 28018 51592 28024
rect 51172 27872 51224 27878
rect 51172 27814 51224 27820
rect 51184 26994 51212 27814
rect 51368 27674 51396 28018
rect 51552 27674 51580 28018
rect 51906 27704 51962 27713
rect 51356 27668 51408 27674
rect 51356 27610 51408 27616
rect 51540 27668 51592 27674
rect 51906 27639 51962 27648
rect 51540 27610 51592 27616
rect 51630 27568 51686 27577
rect 51920 27538 51948 27639
rect 51630 27503 51686 27512
rect 51908 27532 51960 27538
rect 51644 27470 51672 27503
rect 51908 27474 51960 27480
rect 51632 27464 51684 27470
rect 51632 27406 51684 27412
rect 51264 27396 51316 27402
rect 51264 27338 51316 27344
rect 51276 27062 51304 27338
rect 51264 27056 51316 27062
rect 51264 26998 51316 27004
rect 51172 26988 51224 26994
rect 51172 26930 51224 26936
rect 51264 26784 51316 26790
rect 51264 26726 51316 26732
rect 51632 26784 51684 26790
rect 51632 26726 51684 26732
rect 52184 26784 52236 26790
rect 52184 26726 52236 26732
rect 51276 26382 51304 26726
rect 51080 26376 51132 26382
rect 51080 26318 51132 26324
rect 51264 26376 51316 26382
rect 51264 26318 51316 26324
rect 50988 26240 51040 26246
rect 50988 26182 51040 26188
rect 51000 26042 51028 26182
rect 50988 26036 51040 26042
rect 50988 25978 51040 25984
rect 50804 25968 50856 25974
rect 50804 25910 50856 25916
rect 50816 25770 50844 25910
rect 50804 25764 50856 25770
rect 50804 25706 50856 25712
rect 51092 25362 51120 26318
rect 51172 26308 51224 26314
rect 51172 26250 51224 26256
rect 51080 25356 51132 25362
rect 51080 25298 51132 25304
rect 50988 25288 51040 25294
rect 50988 25230 51040 25236
rect 50344 24404 50396 24410
rect 50344 24346 50396 24352
rect 51000 24188 51028 25230
rect 51080 25220 51132 25226
rect 51080 25162 51132 25168
rect 51092 24750 51120 25162
rect 51184 24818 51212 26250
rect 51540 25696 51592 25702
rect 51540 25638 51592 25644
rect 51172 24812 51224 24818
rect 51172 24754 51224 24760
rect 51080 24744 51132 24750
rect 51080 24686 51132 24692
rect 51080 24200 51132 24206
rect 51000 24160 51080 24188
rect 51080 24142 51132 24148
rect 51092 23526 51120 24142
rect 51448 24064 51500 24070
rect 51448 24006 51500 24012
rect 51460 23798 51488 24006
rect 51448 23792 51500 23798
rect 51448 23734 51500 23740
rect 51080 23520 51132 23526
rect 51080 23462 51132 23468
rect 49792 23112 49844 23118
rect 49792 23054 49844 23060
rect 50252 23112 50304 23118
rect 50252 23054 50304 23060
rect 49700 22772 49752 22778
rect 49700 22714 49752 22720
rect 49424 22636 49476 22642
rect 49424 22578 49476 22584
rect 49436 22098 49464 22578
rect 48228 22092 48280 22098
rect 48228 22034 48280 22040
rect 49148 22092 49200 22098
rect 49148 22034 49200 22040
rect 49424 22092 49476 22098
rect 50264 22094 50292 23054
rect 51092 22778 51120 23462
rect 51080 22772 51132 22778
rect 51080 22714 51132 22720
rect 51552 22438 51580 25638
rect 51644 25158 51672 26726
rect 52196 25498 52224 26726
rect 52288 26382 52316 28086
rect 52736 27464 52788 27470
rect 52736 27406 52788 27412
rect 52368 27328 52420 27334
rect 52748 27316 52776 27406
rect 52420 27288 52776 27316
rect 52368 27270 52420 27276
rect 52368 26988 52420 26994
rect 52368 26930 52420 26936
rect 52380 26586 52408 26930
rect 52932 26586 52960 29566
rect 53024 27606 53052 33798
rect 53208 33522 53236 35022
rect 53392 35018 53420 39442
rect 53472 39296 53524 39302
rect 53472 39238 53524 39244
rect 53484 38962 53512 39238
rect 53472 38956 53524 38962
rect 53472 38898 53524 38904
rect 53472 38548 53524 38554
rect 53472 38490 53524 38496
rect 53484 37466 53512 38490
rect 53576 38418 53604 39850
rect 53760 39506 53788 39902
rect 53748 39500 53800 39506
rect 53748 39442 53800 39448
rect 53564 38412 53616 38418
rect 53564 38354 53616 38360
rect 53472 37460 53524 37466
rect 53472 37402 53524 37408
rect 53484 36854 53512 37402
rect 53576 37330 53604 38354
rect 53564 37324 53616 37330
rect 53564 37266 53616 37272
rect 53472 36848 53524 36854
rect 53472 36790 53524 36796
rect 53576 36786 53604 37266
rect 53564 36780 53616 36786
rect 53564 36722 53616 36728
rect 53656 36780 53708 36786
rect 53656 36722 53708 36728
rect 53668 36174 53696 36722
rect 53656 36168 53708 36174
rect 53656 36110 53708 36116
rect 53656 35692 53708 35698
rect 53656 35634 53708 35640
rect 53472 35624 53524 35630
rect 53472 35566 53524 35572
rect 53380 35012 53432 35018
rect 53380 34954 53432 34960
rect 53380 34400 53432 34406
rect 53380 34342 53432 34348
rect 53392 33522 53420 34342
rect 53196 33516 53248 33522
rect 53196 33458 53248 33464
rect 53380 33516 53432 33522
rect 53380 33458 53432 33464
rect 53104 33448 53156 33454
rect 53104 33390 53156 33396
rect 53116 31754 53144 33390
rect 53380 32496 53432 32502
rect 53380 32438 53432 32444
rect 53288 32360 53340 32366
rect 53288 32302 53340 32308
rect 53300 31822 53328 32302
rect 53392 32026 53420 32438
rect 53380 32020 53432 32026
rect 53380 31962 53432 31968
rect 53288 31816 53340 31822
rect 53288 31758 53340 31764
rect 53116 31726 53236 31754
rect 53104 30048 53156 30054
rect 53104 29990 53156 29996
rect 53116 29646 53144 29990
rect 53104 29640 53156 29646
rect 53104 29582 53156 29588
rect 53116 29102 53144 29582
rect 53104 29096 53156 29102
rect 53104 29038 53156 29044
rect 53102 27704 53158 27713
rect 53102 27639 53104 27648
rect 53156 27639 53158 27648
rect 53104 27610 53156 27616
rect 53012 27600 53064 27606
rect 53012 27542 53064 27548
rect 53116 27538 53144 27610
rect 53104 27532 53156 27538
rect 53104 27474 53156 27480
rect 53208 27062 53236 31726
rect 53300 30190 53328 31758
rect 53380 31136 53432 31142
rect 53380 31078 53432 31084
rect 53392 30394 53420 31078
rect 53380 30388 53432 30394
rect 53380 30330 53432 30336
rect 53288 30184 53340 30190
rect 53288 30126 53340 30132
rect 53392 29646 53420 30330
rect 53380 29640 53432 29646
rect 53380 29582 53432 29588
rect 53288 29504 53340 29510
rect 53288 29446 53340 29452
rect 53196 27056 53248 27062
rect 53196 26998 53248 27004
rect 53300 26926 53328 29446
rect 53392 29209 53420 29582
rect 53378 29200 53434 29209
rect 53484 29170 53512 35566
rect 53668 35290 53696 35634
rect 53656 35284 53708 35290
rect 53656 35226 53708 35232
rect 53760 35222 53788 39442
rect 53840 38888 53892 38894
rect 53840 38830 53892 38836
rect 53852 38486 53880 38830
rect 53840 38480 53892 38486
rect 53840 38422 53892 38428
rect 53748 35216 53800 35222
rect 53748 35158 53800 35164
rect 53564 33924 53616 33930
rect 53564 33866 53616 33872
rect 53576 33658 53604 33866
rect 53564 33652 53616 33658
rect 53564 33594 53616 33600
rect 53656 33584 53708 33590
rect 53656 33526 53708 33532
rect 53944 33538 53972 40038
rect 54116 39986 54168 39992
rect 54128 39438 54156 39986
rect 54116 39432 54168 39438
rect 54220 39420 54248 40582
rect 54300 40588 54352 40594
rect 54352 40548 54432 40576
rect 54300 40530 54352 40536
rect 54300 39432 54352 39438
rect 54220 39392 54300 39420
rect 54116 39374 54168 39380
rect 54300 39374 54352 39380
rect 54116 39296 54168 39302
rect 54116 39238 54168 39244
rect 54128 39030 54156 39238
rect 54116 39024 54168 39030
rect 54116 38966 54168 38972
rect 54208 38956 54260 38962
rect 54208 38898 54260 38904
rect 54024 38888 54076 38894
rect 54024 38830 54076 38836
rect 54036 38350 54064 38830
rect 54220 38554 54248 38898
rect 54208 38548 54260 38554
rect 54208 38490 54260 38496
rect 54208 38412 54260 38418
rect 54208 38354 54260 38360
rect 54024 38344 54076 38350
rect 54024 38286 54076 38292
rect 54036 38026 54064 38286
rect 54036 38010 54156 38026
rect 54036 38004 54168 38010
rect 54036 37998 54116 38004
rect 54116 37946 54168 37952
rect 54128 37398 54156 37946
rect 54116 37392 54168 37398
rect 54116 37334 54168 37340
rect 54220 37262 54248 38354
rect 54208 37256 54260 37262
rect 54208 37198 54260 37204
rect 54220 36582 54248 37198
rect 54208 36576 54260 36582
rect 54208 36518 54260 36524
rect 54312 36038 54340 39374
rect 54404 39030 54432 40548
rect 54588 40526 54616 40938
rect 54576 40520 54628 40526
rect 54576 40462 54628 40468
rect 54484 40452 54536 40458
rect 54484 40394 54536 40400
rect 54496 40050 54524 40394
rect 54484 40044 54536 40050
rect 54484 39986 54536 39992
rect 54392 39024 54444 39030
rect 54392 38966 54444 38972
rect 54404 37194 54432 38966
rect 54588 38944 54616 40462
rect 54680 40186 54708 41006
rect 54668 40180 54720 40186
rect 54668 40122 54720 40128
rect 54772 39438 54800 41142
rect 55036 40928 55088 40934
rect 55036 40870 55088 40876
rect 55048 40458 55076 40870
rect 55036 40452 55088 40458
rect 55036 40394 55088 40400
rect 54852 40384 54904 40390
rect 54852 40326 54904 40332
rect 54864 39982 54892 40326
rect 54852 39976 54904 39982
rect 54852 39918 54904 39924
rect 54760 39432 54812 39438
rect 54760 39374 54812 39380
rect 54668 38956 54720 38962
rect 54588 38916 54668 38944
rect 54484 38208 54536 38214
rect 54484 38150 54536 38156
rect 54496 37806 54524 38150
rect 54484 37800 54536 37806
rect 54484 37742 54536 37748
rect 54484 37392 54536 37398
rect 54484 37334 54536 37340
rect 54392 37188 54444 37194
rect 54392 37130 54444 37136
rect 54496 37108 54524 37334
rect 54588 37262 54616 38916
rect 54668 38898 54720 38904
rect 54852 38480 54904 38486
rect 54852 38422 54904 38428
rect 54864 38010 54892 38422
rect 54852 38004 54904 38010
rect 54852 37946 54904 37952
rect 54576 37256 54628 37262
rect 54576 37198 54628 37204
rect 54852 37120 54904 37126
rect 54496 37080 54616 37108
rect 54300 36032 54352 36038
rect 54300 35974 54352 35980
rect 54588 35698 54616 37080
rect 54852 37062 54904 37068
rect 54864 36718 54892 37062
rect 54852 36712 54904 36718
rect 54852 36654 54904 36660
rect 54760 36576 54812 36582
rect 54760 36518 54812 36524
rect 54668 36032 54720 36038
rect 54668 35974 54720 35980
rect 54680 35766 54708 35974
rect 54668 35760 54720 35766
rect 54668 35702 54720 35708
rect 54576 35692 54628 35698
rect 54576 35634 54628 35640
rect 54772 35630 54800 36518
rect 54852 36032 54904 36038
rect 54852 35974 54904 35980
rect 54760 35624 54812 35630
rect 54760 35566 54812 35572
rect 54772 35086 54800 35566
rect 54760 35080 54812 35086
rect 54760 35022 54812 35028
rect 54116 34944 54168 34950
rect 54116 34886 54168 34892
rect 54024 33992 54076 33998
rect 54024 33934 54076 33940
rect 54036 33658 54064 33934
rect 54024 33652 54076 33658
rect 54024 33594 54076 33600
rect 53668 33318 53696 33526
rect 53944 33510 54064 33538
rect 53656 33312 53708 33318
rect 53656 33254 53708 33260
rect 53564 32836 53616 32842
rect 53564 32778 53616 32784
rect 53576 31822 53604 32778
rect 53668 32434 53696 33254
rect 53932 32904 53984 32910
rect 53932 32846 53984 32852
rect 53944 32570 53972 32846
rect 53932 32564 53984 32570
rect 53932 32506 53984 32512
rect 53656 32428 53708 32434
rect 53656 32370 53708 32376
rect 53668 32230 53696 32370
rect 53656 32224 53708 32230
rect 53656 32166 53708 32172
rect 54036 32178 54064 33510
rect 54128 33386 54156 34886
rect 54576 34672 54628 34678
rect 54576 34614 54628 34620
rect 54484 34400 54536 34406
rect 54484 34342 54536 34348
rect 54208 34128 54260 34134
rect 54208 34070 54260 34076
rect 54220 33522 54248 34070
rect 54496 33998 54524 34342
rect 54484 33992 54536 33998
rect 54484 33934 54536 33940
rect 54392 33856 54444 33862
rect 54392 33798 54444 33804
rect 54208 33516 54260 33522
rect 54208 33458 54260 33464
rect 54404 33436 54432 33798
rect 54496 33590 54524 33934
rect 54484 33584 54536 33590
rect 54484 33526 54536 33532
rect 54484 33448 54536 33454
rect 54404 33408 54484 33436
rect 54484 33390 54536 33396
rect 54116 33380 54168 33386
rect 54116 33322 54168 33328
rect 54128 32910 54156 33322
rect 54116 32904 54168 32910
rect 54116 32846 54168 32852
rect 54300 32904 54352 32910
rect 54300 32846 54352 32852
rect 54128 32366 54156 32846
rect 54116 32360 54168 32366
rect 54116 32302 54168 32308
rect 54036 32150 54156 32178
rect 53564 31816 53616 31822
rect 53564 31758 53616 31764
rect 53576 31414 53604 31758
rect 54128 31414 54156 32150
rect 54312 31754 54340 32846
rect 54392 32496 54444 32502
rect 54392 32438 54444 32444
rect 54404 31754 54432 32438
rect 54496 32026 54524 33390
rect 54588 33114 54616 34614
rect 54576 33108 54628 33114
rect 54576 33050 54628 33056
rect 54576 32428 54628 32434
rect 54576 32370 54628 32376
rect 54484 32020 54536 32026
rect 54484 31962 54536 31968
rect 54588 31958 54616 32370
rect 54576 31952 54628 31958
rect 54496 31900 54576 31906
rect 54496 31894 54628 31900
rect 54496 31878 54616 31894
rect 54220 31726 54340 31754
rect 54392 31748 54444 31754
rect 53564 31408 53616 31414
rect 53564 31350 53616 31356
rect 54116 31408 54168 31414
rect 54116 31350 54168 31356
rect 53576 30054 53604 31350
rect 53748 31340 53800 31346
rect 53748 31282 53800 31288
rect 53760 30258 53788 31282
rect 54116 31272 54168 31278
rect 54116 31214 54168 31220
rect 54024 30864 54076 30870
rect 54024 30806 54076 30812
rect 53840 30592 53892 30598
rect 53840 30534 53892 30540
rect 53852 30326 53880 30534
rect 54036 30376 54064 30806
rect 54128 30666 54156 31214
rect 54116 30660 54168 30666
rect 54116 30602 54168 30608
rect 54116 30388 54168 30394
rect 53944 30348 54116 30376
rect 53840 30320 53892 30326
rect 53840 30262 53892 30268
rect 53944 30258 53972 30348
rect 54116 30330 54168 30336
rect 54220 30258 54248 31726
rect 54392 31690 54444 31696
rect 54300 31340 54352 31346
rect 54300 31282 54352 31288
rect 54312 30870 54340 31282
rect 54404 31278 54432 31690
rect 54496 31346 54524 31878
rect 54588 31829 54616 31878
rect 54772 31754 54800 35022
rect 54680 31726 54800 31754
rect 54484 31340 54536 31346
rect 54484 31282 54536 31288
rect 54576 31340 54628 31346
rect 54576 31282 54628 31288
rect 54392 31272 54444 31278
rect 54392 31214 54444 31220
rect 54300 30864 54352 30870
rect 54300 30806 54352 30812
rect 54496 30734 54524 31282
rect 54588 30870 54616 31282
rect 54576 30864 54628 30870
rect 54576 30806 54628 30812
rect 54484 30728 54536 30734
rect 54484 30670 54536 30676
rect 54588 30666 54616 30806
rect 54576 30660 54628 30666
rect 54576 30602 54628 30608
rect 53748 30252 53800 30258
rect 53748 30194 53800 30200
rect 53932 30252 53984 30258
rect 53932 30194 53984 30200
rect 54208 30252 54260 30258
rect 54208 30194 54260 30200
rect 53564 30048 53616 30054
rect 53564 29990 53616 29996
rect 53760 29850 53788 30194
rect 53748 29844 53800 29850
rect 53748 29786 53800 29792
rect 53564 29708 53616 29714
rect 53564 29650 53616 29656
rect 53576 29578 53604 29650
rect 53564 29572 53616 29578
rect 53564 29514 53616 29520
rect 53378 29135 53434 29144
rect 53472 29164 53524 29170
rect 54392 29164 54444 29170
rect 53524 29124 53604 29152
rect 53472 29106 53524 29112
rect 53472 28960 53524 28966
rect 53472 28902 53524 28908
rect 53484 28558 53512 28902
rect 53380 28552 53432 28558
rect 53380 28494 53432 28500
rect 53472 28552 53524 28558
rect 53472 28494 53524 28500
rect 53392 28218 53420 28494
rect 53380 28212 53432 28218
rect 53380 28154 53432 28160
rect 53576 28150 53604 29124
rect 54392 29106 54444 29112
rect 53656 28960 53708 28966
rect 53656 28902 53708 28908
rect 53668 28558 53696 28902
rect 54404 28694 54432 29106
rect 54392 28688 54444 28694
rect 54392 28630 54444 28636
rect 53656 28552 53708 28558
rect 53656 28494 53708 28500
rect 54116 28552 54168 28558
rect 54116 28494 54168 28500
rect 54024 28484 54076 28490
rect 54024 28426 54076 28432
rect 53932 28416 53984 28422
rect 53932 28358 53984 28364
rect 53564 28144 53616 28150
rect 53564 28086 53616 28092
rect 53472 27532 53524 27538
rect 53472 27474 53524 27480
rect 53288 26920 53340 26926
rect 53288 26862 53340 26868
rect 53484 26790 53512 27474
rect 53576 26994 53604 28086
rect 53944 27470 53972 28358
rect 54036 28150 54064 28426
rect 54024 28144 54076 28150
rect 54024 28086 54076 28092
rect 54128 27946 54156 28494
rect 54404 28082 54432 28630
rect 54588 28370 54616 30602
rect 54680 29714 54708 31726
rect 54760 31136 54812 31142
rect 54760 31078 54812 31084
rect 54772 30734 54800 31078
rect 54760 30728 54812 30734
rect 54760 30670 54812 30676
rect 54668 29708 54720 29714
rect 54668 29650 54720 29656
rect 54680 29238 54708 29650
rect 54668 29232 54720 29238
rect 54668 29174 54720 29180
rect 54496 28342 54616 28370
rect 54392 28076 54444 28082
rect 54392 28018 54444 28024
rect 54116 27940 54168 27946
rect 54116 27882 54168 27888
rect 53932 27464 53984 27470
rect 53932 27406 53984 27412
rect 54300 27464 54352 27470
rect 54300 27406 54352 27412
rect 53564 26988 53616 26994
rect 53564 26930 53616 26936
rect 54312 26858 54340 27406
rect 54496 27130 54524 28342
rect 54680 28200 54708 29174
rect 54864 29050 54892 35974
rect 54944 33448 54996 33454
rect 54944 33390 54996 33396
rect 54956 32502 54984 33390
rect 54944 32496 54996 32502
rect 54944 32438 54996 32444
rect 54956 31822 54984 32438
rect 54944 31816 54996 31822
rect 54944 31758 54996 31764
rect 54956 30784 54984 31758
rect 55048 31686 55076 40394
rect 55220 38752 55272 38758
rect 55220 38694 55272 38700
rect 55232 38418 55260 38694
rect 55312 38548 55364 38554
rect 55312 38490 55364 38496
rect 55220 38412 55272 38418
rect 55220 38354 55272 38360
rect 55128 36576 55180 36582
rect 55128 36518 55180 36524
rect 55140 36174 55168 36518
rect 55128 36168 55180 36174
rect 55128 36110 55180 36116
rect 55220 36032 55272 36038
rect 55220 35974 55272 35980
rect 55036 31680 55088 31686
rect 55036 31622 55088 31628
rect 55048 31346 55076 31622
rect 55036 31340 55088 31346
rect 55036 31282 55088 31288
rect 54956 30756 55076 30784
rect 54944 30660 54996 30666
rect 54944 30602 54996 30608
rect 54956 30258 54984 30602
rect 55048 30326 55076 30756
rect 55036 30320 55088 30326
rect 55036 30262 55088 30268
rect 54944 30252 54996 30258
rect 54944 30194 54996 30200
rect 55128 30048 55180 30054
rect 55128 29990 55180 29996
rect 55140 29714 55168 29990
rect 55128 29708 55180 29714
rect 55128 29650 55180 29656
rect 55232 29306 55260 35974
rect 55324 30326 55352 38490
rect 55404 35488 55456 35494
rect 55404 35430 55456 35436
rect 55416 34490 55444 35430
rect 55508 35154 55536 43794
rect 55784 43790 55812 44338
rect 56140 44328 56192 44334
rect 56140 44270 56192 44276
rect 55772 43784 55824 43790
rect 55772 43726 55824 43732
rect 55588 41064 55640 41070
rect 55588 41006 55640 41012
rect 55600 40526 55628 41006
rect 55588 40520 55640 40526
rect 55588 40462 55640 40468
rect 55680 40112 55732 40118
rect 55680 40054 55732 40060
rect 55588 39840 55640 39846
rect 55588 39782 55640 39788
rect 55600 39370 55628 39782
rect 55588 39364 55640 39370
rect 55588 39306 55640 39312
rect 55600 38554 55628 39306
rect 55588 38548 55640 38554
rect 55588 38490 55640 38496
rect 55692 38350 55720 40054
rect 55956 39500 56008 39506
rect 55956 39442 56008 39448
rect 55772 39432 55824 39438
rect 55772 39374 55824 39380
rect 55784 39098 55812 39374
rect 55772 39092 55824 39098
rect 55772 39034 55824 39040
rect 55680 38344 55732 38350
rect 55680 38286 55732 38292
rect 55784 37262 55812 39034
rect 55968 37874 55996 39442
rect 56048 39296 56100 39302
rect 56048 39238 56100 39244
rect 56060 38894 56088 39238
rect 56048 38888 56100 38894
rect 56048 38830 56100 38836
rect 56048 38208 56100 38214
rect 56048 38150 56100 38156
rect 55956 37868 56008 37874
rect 55956 37810 56008 37816
rect 56060 37806 56088 38150
rect 56152 38026 56180 44270
rect 57244 42696 57296 42702
rect 57244 42638 57296 42644
rect 56692 42560 56744 42566
rect 56692 42502 56744 42508
rect 57060 42560 57112 42566
rect 57060 42502 57112 42508
rect 56232 41608 56284 41614
rect 56232 41550 56284 41556
rect 56244 41274 56272 41550
rect 56232 41268 56284 41274
rect 56232 41210 56284 41216
rect 56600 40452 56652 40458
rect 56600 40394 56652 40400
rect 56612 40050 56640 40394
rect 56600 40044 56652 40050
rect 56600 39986 56652 39992
rect 56508 39296 56560 39302
rect 56508 39238 56560 39244
rect 56520 38962 56548 39238
rect 56508 38956 56560 38962
rect 56508 38898 56560 38904
rect 56152 37998 56272 38026
rect 56140 37936 56192 37942
rect 56140 37878 56192 37884
rect 55864 37800 55916 37806
rect 55864 37742 55916 37748
rect 56048 37800 56100 37806
rect 56048 37742 56100 37748
rect 55876 37330 55904 37742
rect 55864 37324 55916 37330
rect 55864 37266 55916 37272
rect 55772 37256 55824 37262
rect 55772 37198 55824 37204
rect 56152 36174 56180 37878
rect 56244 36802 56272 37998
rect 56324 37868 56376 37874
rect 56324 37810 56376 37816
rect 56336 37466 56364 37810
rect 56324 37460 56376 37466
rect 56324 37402 56376 37408
rect 56244 36774 56364 36802
rect 56232 36644 56284 36650
rect 56232 36586 56284 36592
rect 56140 36168 56192 36174
rect 56140 36110 56192 36116
rect 56152 35698 56180 36110
rect 56140 35692 56192 35698
rect 56140 35634 56192 35640
rect 55772 35216 55824 35222
rect 55772 35158 55824 35164
rect 55496 35148 55548 35154
rect 55496 35090 55548 35096
rect 55508 34610 55536 35090
rect 55784 35086 55812 35158
rect 55772 35080 55824 35086
rect 55772 35022 55824 35028
rect 56140 35080 56192 35086
rect 56140 35022 56192 35028
rect 55496 34604 55548 34610
rect 55496 34546 55548 34552
rect 55588 34536 55640 34542
rect 55416 34462 55536 34490
rect 55588 34478 55640 34484
rect 55404 33380 55456 33386
rect 55404 33322 55456 33328
rect 55416 31890 55444 33322
rect 55404 31884 55456 31890
rect 55404 31826 55456 31832
rect 55312 30320 55364 30326
rect 55312 30262 55364 30268
rect 55508 30190 55536 34462
rect 55600 33114 55628 34478
rect 55784 33930 55812 35022
rect 55956 34944 56008 34950
rect 55956 34886 56008 34892
rect 55968 33998 55996 34886
rect 56152 34542 56180 35022
rect 56140 34536 56192 34542
rect 56140 34478 56192 34484
rect 56048 34400 56100 34406
rect 56048 34342 56100 34348
rect 56060 33998 56088 34342
rect 56244 33998 56272 36586
rect 56336 35086 56364 36774
rect 56600 36576 56652 36582
rect 56600 36518 56652 36524
rect 56612 35222 56640 36518
rect 56704 35766 56732 42502
rect 56876 39432 56928 39438
rect 56876 39374 56928 39380
rect 56888 39098 56916 39374
rect 56876 39092 56928 39098
rect 56876 39034 56928 39040
rect 56876 36032 56928 36038
rect 56876 35974 56928 35980
rect 56692 35760 56744 35766
rect 56692 35702 56744 35708
rect 56600 35216 56652 35222
rect 56600 35158 56652 35164
rect 56324 35080 56376 35086
rect 56324 35022 56376 35028
rect 56336 34746 56364 35022
rect 56324 34740 56376 34746
rect 56324 34682 56376 34688
rect 56336 34610 56364 34682
rect 56324 34604 56376 34610
rect 56324 34546 56376 34552
rect 55956 33992 56008 33998
rect 55956 33934 56008 33940
rect 56048 33992 56100 33998
rect 56048 33934 56100 33940
rect 56232 33992 56284 33998
rect 56232 33934 56284 33940
rect 56612 33930 56640 35158
rect 55772 33924 55824 33930
rect 55772 33866 55824 33872
rect 55864 33924 55916 33930
rect 55864 33866 55916 33872
rect 56600 33924 56652 33930
rect 56600 33866 56652 33872
rect 55588 33108 55640 33114
rect 55588 33050 55640 33056
rect 55772 33040 55824 33046
rect 55772 32982 55824 32988
rect 55784 32910 55812 32982
rect 55772 32904 55824 32910
rect 55772 32846 55824 32852
rect 55784 32502 55812 32846
rect 55772 32496 55824 32502
rect 55772 32438 55824 32444
rect 55588 32428 55640 32434
rect 55588 32370 55640 32376
rect 55600 31822 55628 32370
rect 55588 31816 55640 31822
rect 55588 31758 55640 31764
rect 55600 31278 55628 31758
rect 55588 31272 55640 31278
rect 55588 31214 55640 31220
rect 55496 30184 55548 30190
rect 55496 30126 55548 30132
rect 55600 30036 55628 31214
rect 55876 30938 55904 33866
rect 56612 33522 56640 33866
rect 56600 33516 56652 33522
rect 56600 33458 56652 33464
rect 56232 32904 56284 32910
rect 56232 32846 56284 32852
rect 56244 32570 56272 32846
rect 56232 32564 56284 32570
rect 56232 32506 56284 32512
rect 56324 32496 56376 32502
rect 56612 32450 56640 33458
rect 56704 33386 56732 35702
rect 56784 33856 56836 33862
rect 56784 33798 56836 33804
rect 56796 33454 56824 33798
rect 56784 33448 56836 33454
rect 56784 33390 56836 33396
rect 56692 33380 56744 33386
rect 56692 33322 56744 33328
rect 56704 33114 56732 33322
rect 56692 33108 56744 33114
rect 56692 33050 56744 33056
rect 56784 32972 56836 32978
rect 56784 32914 56836 32920
rect 56324 32438 56376 32444
rect 55956 32428 56008 32434
rect 55956 32370 56008 32376
rect 55968 32298 55996 32370
rect 55956 32292 56008 32298
rect 55956 32234 56008 32240
rect 55968 31822 55996 32234
rect 56336 31890 56364 32438
rect 56416 32428 56468 32434
rect 56416 32370 56468 32376
rect 56520 32422 56640 32450
rect 56796 32434 56824 32914
rect 56784 32428 56836 32434
rect 56428 32026 56456 32370
rect 56520 32178 56548 32422
rect 56784 32370 56836 32376
rect 56520 32150 56732 32178
rect 56416 32020 56468 32026
rect 56416 31962 56468 31968
rect 56324 31884 56376 31890
rect 56324 31826 56376 31832
rect 55956 31816 56008 31822
rect 55956 31758 56008 31764
rect 56140 31816 56192 31822
rect 56140 31758 56192 31764
rect 56152 31346 56180 31758
rect 56336 31414 56364 31826
rect 56324 31408 56376 31414
rect 56324 31350 56376 31356
rect 56140 31340 56192 31346
rect 56140 31282 56192 31288
rect 55864 30932 55916 30938
rect 55864 30874 55916 30880
rect 56152 30258 56180 31282
rect 55772 30252 55824 30258
rect 55772 30194 55824 30200
rect 56140 30252 56192 30258
rect 56140 30194 56192 30200
rect 55324 30008 55628 30036
rect 55324 29578 55352 30008
rect 55784 29730 55812 30194
rect 56048 30116 56100 30122
rect 56048 30058 56100 30064
rect 55956 30048 56008 30054
rect 55956 29990 56008 29996
rect 55508 29702 55812 29730
rect 55508 29646 55536 29702
rect 55784 29646 55812 29702
rect 55496 29640 55548 29646
rect 55496 29582 55548 29588
rect 55588 29640 55640 29646
rect 55588 29582 55640 29588
rect 55772 29640 55824 29646
rect 55772 29582 55824 29588
rect 55312 29572 55364 29578
rect 55312 29514 55364 29520
rect 55496 29504 55548 29510
rect 55496 29446 55548 29452
rect 55220 29300 55272 29306
rect 55220 29242 55272 29248
rect 54772 29022 54892 29050
rect 54772 28558 54800 29022
rect 54852 28960 54904 28966
rect 54852 28902 54904 28908
rect 54864 28626 54892 28902
rect 54852 28620 54904 28626
rect 54852 28562 54904 28568
rect 54760 28552 54812 28558
rect 54760 28494 54812 28500
rect 54588 28172 54708 28200
rect 54484 27124 54536 27130
rect 54484 27066 54536 27072
rect 54300 26852 54352 26858
rect 54300 26794 54352 26800
rect 53472 26784 53524 26790
rect 53472 26726 53524 26732
rect 53564 26784 53616 26790
rect 53564 26726 53616 26732
rect 53576 26586 53604 26726
rect 54312 26586 54340 26794
rect 52368 26580 52420 26586
rect 52368 26522 52420 26528
rect 52920 26580 52972 26586
rect 52920 26522 52972 26528
rect 53564 26580 53616 26586
rect 53564 26522 53616 26528
rect 54300 26580 54352 26586
rect 54300 26522 54352 26528
rect 52276 26376 52328 26382
rect 52276 26318 52328 26324
rect 52380 26042 52408 26522
rect 54496 26518 54524 27066
rect 54484 26512 54536 26518
rect 54484 26454 54536 26460
rect 54588 26042 54616 28172
rect 54772 27452 54800 28494
rect 55232 28218 55260 29242
rect 55402 29200 55458 29209
rect 55508 29170 55536 29446
rect 55600 29238 55628 29582
rect 55588 29232 55640 29238
rect 55588 29174 55640 29180
rect 55968 29170 55996 29990
rect 56060 29646 56088 30058
rect 56048 29640 56100 29646
rect 56048 29582 56100 29588
rect 55402 29135 55404 29144
rect 55456 29135 55458 29144
rect 55496 29164 55548 29170
rect 55404 29106 55456 29112
rect 55496 29106 55548 29112
rect 55956 29164 56008 29170
rect 56060 29152 56088 29582
rect 56140 29164 56192 29170
rect 56060 29124 56140 29152
rect 55956 29106 56008 29112
rect 56140 29106 56192 29112
rect 55588 28960 55640 28966
rect 55588 28902 55640 28908
rect 55220 28212 55272 28218
rect 55220 28154 55272 28160
rect 55600 28014 55628 28902
rect 55588 28008 55640 28014
rect 55588 27950 55640 27956
rect 55864 27872 55916 27878
rect 55864 27814 55916 27820
rect 55876 27470 55904 27814
rect 54852 27464 54904 27470
rect 54772 27424 54852 27452
rect 54852 27406 54904 27412
rect 55864 27464 55916 27470
rect 55864 27406 55916 27412
rect 54760 27328 54812 27334
rect 54760 27270 54812 27276
rect 54772 27130 54800 27270
rect 54760 27124 54812 27130
rect 54760 27066 54812 27072
rect 54668 26988 54720 26994
rect 54668 26930 54720 26936
rect 54680 26586 54708 26930
rect 54668 26580 54720 26586
rect 54668 26522 54720 26528
rect 54864 26450 54892 27406
rect 55036 27328 55088 27334
rect 55036 27270 55088 27276
rect 55128 27328 55180 27334
rect 55128 27270 55180 27276
rect 55048 27062 55076 27270
rect 55140 27062 55168 27270
rect 55876 27062 55904 27406
rect 55036 27056 55088 27062
rect 55036 26998 55088 27004
rect 55128 27056 55180 27062
rect 55128 26998 55180 27004
rect 55864 27056 55916 27062
rect 55864 26998 55916 27004
rect 54852 26444 54904 26450
rect 54852 26386 54904 26392
rect 56152 26042 56180 29106
rect 56336 27878 56364 31350
rect 56508 30660 56560 30666
rect 56508 30602 56560 30608
rect 56416 30184 56468 30190
rect 56416 30126 56468 30132
rect 56428 29578 56456 30126
rect 56520 29782 56548 30602
rect 56600 30320 56652 30326
rect 56600 30262 56652 30268
rect 56508 29776 56560 29782
rect 56508 29718 56560 29724
rect 56416 29572 56468 29578
rect 56416 29514 56468 29520
rect 56324 27872 56376 27878
rect 56324 27814 56376 27820
rect 56336 26586 56364 27814
rect 56520 27470 56548 29718
rect 56612 28422 56640 30262
rect 56704 29238 56732 32150
rect 56796 31414 56824 32370
rect 56784 31408 56836 31414
rect 56784 31350 56836 31356
rect 56888 29782 56916 35974
rect 56968 34944 57020 34950
rect 56968 34886 57020 34892
rect 56980 33998 57008 34886
rect 57072 34542 57100 42502
rect 57256 41682 57284 42638
rect 57336 42356 57388 42362
rect 57336 42298 57388 42304
rect 57244 41676 57296 41682
rect 57244 41618 57296 41624
rect 57244 40520 57296 40526
rect 57244 40462 57296 40468
rect 57256 40186 57284 40462
rect 57244 40180 57296 40186
rect 57244 40122 57296 40128
rect 57244 40044 57296 40050
rect 57244 39986 57296 39992
rect 57256 39438 57284 39986
rect 57244 39432 57296 39438
rect 57244 39374 57296 39380
rect 57244 37664 57296 37670
rect 57244 37606 57296 37612
rect 57152 35080 57204 35086
rect 57152 35022 57204 35028
rect 57164 34746 57192 35022
rect 57152 34740 57204 34746
rect 57152 34682 57204 34688
rect 57060 34536 57112 34542
rect 57060 34478 57112 34484
rect 56968 33992 57020 33998
rect 56968 33934 57020 33940
rect 57072 33658 57100 34478
rect 57060 33652 57112 33658
rect 57060 33594 57112 33600
rect 57152 32972 57204 32978
rect 57152 32914 57204 32920
rect 57060 32836 57112 32842
rect 57060 32778 57112 32784
rect 57072 32434 57100 32778
rect 57164 32570 57192 32914
rect 57152 32564 57204 32570
rect 57152 32506 57204 32512
rect 57060 32428 57112 32434
rect 57060 32370 57112 32376
rect 57072 31414 57100 32370
rect 57060 31408 57112 31414
rect 57060 31350 57112 31356
rect 57152 31136 57204 31142
rect 57152 31078 57204 31084
rect 57164 30734 57192 31078
rect 57152 30728 57204 30734
rect 57152 30670 57204 30676
rect 57060 30592 57112 30598
rect 57060 30534 57112 30540
rect 57072 30190 57100 30534
rect 57060 30184 57112 30190
rect 57060 30126 57112 30132
rect 57256 29866 57284 37606
rect 57348 35766 57376 42298
rect 57428 41676 57480 41682
rect 57428 41618 57480 41624
rect 57440 40526 57468 41618
rect 57428 40520 57480 40526
rect 57428 40462 57480 40468
rect 58256 40384 58308 40390
rect 58256 40326 58308 40332
rect 57704 37732 57756 37738
rect 57704 37674 57756 37680
rect 57716 36174 57744 37674
rect 57980 37120 58032 37126
rect 57980 37062 58032 37068
rect 57992 36582 58020 37062
rect 57980 36576 58032 36582
rect 57980 36518 58032 36524
rect 57428 36168 57480 36174
rect 57428 36110 57480 36116
rect 57704 36168 57756 36174
rect 57704 36110 57756 36116
rect 57440 35834 57468 36110
rect 57428 35828 57480 35834
rect 57428 35770 57480 35776
rect 57336 35760 57388 35766
rect 57336 35702 57388 35708
rect 57348 35170 57376 35702
rect 57704 35488 57756 35494
rect 57704 35430 57756 35436
rect 57348 35142 57468 35170
rect 57336 35080 57388 35086
rect 57336 35022 57388 35028
rect 57348 34406 57376 35022
rect 57336 34400 57388 34406
rect 57336 34342 57388 34348
rect 57440 33810 57468 35142
rect 57716 35018 57744 35430
rect 58072 35216 58124 35222
rect 58072 35158 58124 35164
rect 57980 35148 58032 35154
rect 57980 35090 58032 35096
rect 57704 35012 57756 35018
rect 57704 34954 57756 34960
rect 57716 34202 57744 34954
rect 57992 34678 58020 35090
rect 57980 34672 58032 34678
rect 57980 34614 58032 34620
rect 58084 34610 58112 35158
rect 58072 34604 58124 34610
rect 58072 34546 58124 34552
rect 57704 34196 57756 34202
rect 57704 34138 57756 34144
rect 57348 33782 57468 33810
rect 57348 32502 57376 33782
rect 57428 33652 57480 33658
rect 57428 33594 57480 33600
rect 57440 32910 57468 33594
rect 57520 33516 57572 33522
rect 57520 33458 57572 33464
rect 57532 33114 57560 33458
rect 57520 33108 57572 33114
rect 57520 33050 57572 33056
rect 57428 32904 57480 32910
rect 57428 32846 57480 32852
rect 57336 32496 57388 32502
rect 57336 32438 57388 32444
rect 57612 31816 57664 31822
rect 57612 31758 57664 31764
rect 57624 31210 57652 31758
rect 57716 31754 57744 34138
rect 57888 33448 57940 33454
rect 57980 33448 58032 33454
rect 57940 33408 57980 33436
rect 57888 33390 57940 33396
rect 57980 33390 58032 33396
rect 57980 33312 58032 33318
rect 57980 33254 58032 33260
rect 57992 32978 58020 33254
rect 57980 32972 58032 32978
rect 57980 32914 58032 32920
rect 58268 32842 58296 40326
rect 58440 39296 58492 39302
rect 58440 39238 58492 39244
rect 58256 32836 58308 32842
rect 58256 32778 58308 32784
rect 58164 32768 58216 32774
rect 58164 32710 58216 32716
rect 57980 32224 58032 32230
rect 57980 32166 58032 32172
rect 57716 31748 57848 31754
rect 57716 31726 57796 31748
rect 57796 31690 57848 31696
rect 57992 31686 58020 32166
rect 58072 31952 58124 31958
rect 58072 31894 58124 31900
rect 57980 31680 58032 31686
rect 57980 31622 58032 31628
rect 58084 31278 58112 31894
rect 57888 31272 57940 31278
rect 57888 31214 57940 31220
rect 58072 31272 58124 31278
rect 58072 31214 58124 31220
rect 57612 31204 57664 31210
rect 57612 31146 57664 31152
rect 57624 30938 57652 31146
rect 57796 31136 57848 31142
rect 57796 31078 57848 31084
rect 57612 30932 57664 30938
rect 57612 30874 57664 30880
rect 57336 30796 57388 30802
rect 57336 30738 57388 30744
rect 57348 30258 57376 30738
rect 57336 30252 57388 30258
rect 57336 30194 57388 30200
rect 57520 30116 57572 30122
rect 57520 30058 57572 30064
rect 57164 29838 57284 29866
rect 56876 29776 56928 29782
rect 56876 29718 56928 29724
rect 56692 29232 56744 29238
rect 56692 29174 56744 29180
rect 56600 28416 56652 28422
rect 56600 28358 56652 28364
rect 56508 27464 56560 27470
rect 56508 27406 56560 27412
rect 56612 26790 56640 28358
rect 56888 27402 56916 29718
rect 57164 28082 57192 29838
rect 57244 29708 57296 29714
rect 57244 29650 57296 29656
rect 57256 28558 57284 29650
rect 57336 29164 57388 29170
rect 57336 29106 57388 29112
rect 57348 28694 57376 29106
rect 57336 28688 57388 28694
rect 57336 28630 57388 28636
rect 57244 28552 57296 28558
rect 57244 28494 57296 28500
rect 57244 28416 57296 28422
rect 57244 28358 57296 28364
rect 57152 28076 57204 28082
rect 57152 28018 57204 28024
rect 57256 28014 57284 28358
rect 57244 28008 57296 28014
rect 57244 27950 57296 27956
rect 57348 27946 57376 28630
rect 57532 28626 57560 30058
rect 57520 28620 57572 28626
rect 57520 28562 57572 28568
rect 57336 27940 57388 27946
rect 57336 27882 57388 27888
rect 57704 27872 57756 27878
rect 57704 27814 57756 27820
rect 57716 27538 57744 27814
rect 57808 27606 57836 31078
rect 57900 30394 57928 31214
rect 57888 30388 57940 30394
rect 57888 30330 57940 30336
rect 57796 27600 57848 27606
rect 57796 27542 57848 27548
rect 57704 27532 57756 27538
rect 57704 27474 57756 27480
rect 56876 27396 56928 27402
rect 56876 27338 56928 27344
rect 56888 27130 56916 27338
rect 56876 27124 56928 27130
rect 56876 27066 56928 27072
rect 57900 27062 57928 30330
rect 57980 29640 58032 29646
rect 57980 29582 58032 29588
rect 56692 27056 56744 27062
rect 56692 26998 56744 27004
rect 57888 27056 57940 27062
rect 57888 26998 57940 27004
rect 56600 26784 56652 26790
rect 56600 26726 56652 26732
rect 56704 26586 56732 26998
rect 56324 26580 56376 26586
rect 56324 26522 56376 26528
rect 56692 26580 56744 26586
rect 56692 26522 56744 26528
rect 52368 26036 52420 26042
rect 52368 25978 52420 25984
rect 54576 26036 54628 26042
rect 54576 25978 54628 25984
rect 56140 26036 56192 26042
rect 56140 25978 56192 25984
rect 52184 25492 52236 25498
rect 52184 25434 52236 25440
rect 57992 25430 58020 29582
rect 58072 28008 58124 28014
rect 58072 27950 58124 27956
rect 58084 27674 58112 27950
rect 58072 27668 58124 27674
rect 58072 27610 58124 27616
rect 58072 27464 58124 27470
rect 58072 27406 58124 27412
rect 58084 26790 58112 27406
rect 58176 27402 58204 32710
rect 58268 31822 58296 32778
rect 58348 31884 58400 31890
rect 58348 31826 58400 31832
rect 58256 31816 58308 31822
rect 58256 31758 58308 31764
rect 58256 29504 58308 29510
rect 58256 29446 58308 29452
rect 58268 29345 58296 29446
rect 58254 29336 58310 29345
rect 58360 29306 58388 31826
rect 58452 30802 58480 39238
rect 58532 31816 58584 31822
rect 58532 31758 58584 31764
rect 58544 31346 58572 31758
rect 58532 31340 58584 31346
rect 58532 31282 58584 31288
rect 58636 31249 58664 56646
rect 58622 31240 58678 31249
rect 58622 31175 58678 31184
rect 58440 30796 58492 30802
rect 58440 30738 58492 30744
rect 58254 29271 58310 29280
rect 58348 29300 58400 29306
rect 58348 29242 58400 29248
rect 58348 28076 58400 28082
rect 58348 28018 58400 28024
rect 58360 27470 58388 28018
rect 58348 27464 58400 27470
rect 58348 27406 58400 27412
rect 58164 27396 58216 27402
rect 58164 27338 58216 27344
rect 58256 27328 58308 27334
rect 58256 27270 58308 27276
rect 58072 26784 58124 26790
rect 58072 26726 58124 26732
rect 58084 26314 58112 26726
rect 58072 26308 58124 26314
rect 58072 26250 58124 26256
rect 58268 26042 58296 27270
rect 58256 26036 58308 26042
rect 58256 25978 58308 25984
rect 52644 25424 52696 25430
rect 52644 25366 52696 25372
rect 57980 25424 58032 25430
rect 57980 25366 58032 25372
rect 51816 25288 51868 25294
rect 51816 25230 51868 25236
rect 51632 25152 51684 25158
rect 51632 25094 51684 25100
rect 51644 24750 51672 25094
rect 51632 24744 51684 24750
rect 51632 24686 51684 24692
rect 51828 23730 51856 25230
rect 52656 24818 52684 25366
rect 52644 24812 52696 24818
rect 52644 24754 52696 24760
rect 51816 23724 51868 23730
rect 51816 23666 51868 23672
rect 51828 23322 51856 23666
rect 51816 23316 51868 23322
rect 51816 23258 51868 23264
rect 51540 22432 51592 22438
rect 51540 22374 51592 22380
rect 58164 22432 58216 22438
rect 58164 22374 58216 22380
rect 50264 22066 50384 22094
rect 49424 22034 49476 22040
rect 47768 21684 47820 21690
rect 47768 21626 47820 21632
rect 47308 21140 47360 21146
rect 47308 21082 47360 21088
rect 50356 20942 50384 22066
rect 50344 20936 50396 20942
rect 50344 20878 50396 20884
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34716 6886 34836 6914
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 34716 2650 34744 6886
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 58176 2650 58204 22374
rect 58624 2848 58676 2854
rect 58624 2790 58676 2796
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 34704 2644 34756 2650
rect 34704 2586 34756 2592
rect 58164 2644 58216 2650
rect 58164 2586 58216 2592
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 1596 1358 1624 2382
rect 58636 2378 58664 2790
rect 58624 2372 58676 2378
rect 58624 2314 58676 2320
rect 29000 2304 29052 2310
rect 29000 2246 29052 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 20 1352 72 1358
rect 20 1294 72 1300
rect 1584 1352 1636 1358
rect 1584 1294 1636 1300
rect 32 800 60 1294
rect 29012 800 29040 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 58636 800 58664 2314
rect 18 200 74 800
rect 28998 200 29054 800
rect 58622 200 58678 800
<< via2 >>
rect 4880 57690 4936 57692
rect 4960 57690 5016 57692
rect 5040 57690 5096 57692
rect 5120 57690 5176 57692
rect 4880 57638 4926 57690
rect 4926 57638 4936 57690
rect 4960 57638 4990 57690
rect 4990 57638 5002 57690
rect 5002 57638 5016 57690
rect 5040 57638 5054 57690
rect 5054 57638 5066 57690
rect 5066 57638 5096 57690
rect 5120 57638 5130 57690
rect 5130 57638 5176 57690
rect 4880 57636 4936 57638
rect 4960 57636 5016 57638
rect 5040 57636 5096 57638
rect 5120 57636 5176 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4880 56602 4936 56604
rect 4960 56602 5016 56604
rect 5040 56602 5096 56604
rect 5120 56602 5176 56604
rect 4880 56550 4926 56602
rect 4926 56550 4936 56602
rect 4960 56550 4990 56602
rect 4990 56550 5002 56602
rect 5002 56550 5016 56602
rect 5040 56550 5054 56602
rect 5054 56550 5066 56602
rect 5066 56550 5096 56602
rect 5120 56550 5130 56602
rect 5130 56550 5176 56602
rect 4880 56548 4936 56550
rect 4960 56548 5016 56550
rect 5040 56548 5096 56550
rect 5120 56548 5176 56550
rect 35600 57690 35656 57692
rect 35680 57690 35736 57692
rect 35760 57690 35816 57692
rect 35840 57690 35896 57692
rect 35600 57638 35646 57690
rect 35646 57638 35656 57690
rect 35680 57638 35710 57690
rect 35710 57638 35722 57690
rect 35722 57638 35736 57690
rect 35760 57638 35774 57690
rect 35774 57638 35786 57690
rect 35786 57638 35816 57690
rect 35840 57638 35850 57690
rect 35850 57638 35896 57690
rect 35600 57636 35656 57638
rect 35680 57636 35736 57638
rect 35760 57636 35816 57638
rect 35840 57636 35896 57638
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 35600 56602 35656 56604
rect 35680 56602 35736 56604
rect 35760 56602 35816 56604
rect 35840 56602 35896 56604
rect 35600 56550 35646 56602
rect 35646 56550 35656 56602
rect 35680 56550 35710 56602
rect 35710 56550 35722 56602
rect 35722 56550 35736 56602
rect 35760 56550 35774 56602
rect 35774 56550 35786 56602
rect 35786 56550 35816 56602
rect 35840 56550 35850 56602
rect 35850 56550 35896 56602
rect 35600 56548 35656 56550
rect 35680 56548 35736 56550
rect 35760 56548 35816 56550
rect 35840 56548 35896 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4880 55514 4936 55516
rect 4960 55514 5016 55516
rect 5040 55514 5096 55516
rect 5120 55514 5176 55516
rect 4880 55462 4926 55514
rect 4926 55462 4936 55514
rect 4960 55462 4990 55514
rect 4990 55462 5002 55514
rect 5002 55462 5016 55514
rect 5040 55462 5054 55514
rect 5054 55462 5066 55514
rect 5066 55462 5096 55514
rect 5120 55462 5130 55514
rect 5130 55462 5176 55514
rect 4880 55460 4936 55462
rect 4960 55460 5016 55462
rect 5040 55460 5096 55462
rect 5120 55460 5176 55462
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 35600 55514 35656 55516
rect 35680 55514 35736 55516
rect 35760 55514 35816 55516
rect 35840 55514 35896 55516
rect 35600 55462 35646 55514
rect 35646 55462 35656 55514
rect 35680 55462 35710 55514
rect 35710 55462 35722 55514
rect 35722 55462 35736 55514
rect 35760 55462 35774 55514
rect 35774 55462 35786 55514
rect 35786 55462 35816 55514
rect 35840 55462 35850 55514
rect 35850 55462 35896 55514
rect 35600 55460 35656 55462
rect 35680 55460 35736 55462
rect 35760 55460 35816 55462
rect 35840 55460 35896 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4880 54426 4936 54428
rect 4960 54426 5016 54428
rect 5040 54426 5096 54428
rect 5120 54426 5176 54428
rect 4880 54374 4926 54426
rect 4926 54374 4936 54426
rect 4960 54374 4990 54426
rect 4990 54374 5002 54426
rect 5002 54374 5016 54426
rect 5040 54374 5054 54426
rect 5054 54374 5066 54426
rect 5066 54374 5096 54426
rect 5120 54374 5130 54426
rect 5130 54374 5176 54426
rect 4880 54372 4936 54374
rect 4960 54372 5016 54374
rect 5040 54372 5096 54374
rect 5120 54372 5176 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4880 53338 4936 53340
rect 4960 53338 5016 53340
rect 5040 53338 5096 53340
rect 5120 53338 5176 53340
rect 4880 53286 4926 53338
rect 4926 53286 4936 53338
rect 4960 53286 4990 53338
rect 4990 53286 5002 53338
rect 5002 53286 5016 53338
rect 5040 53286 5054 53338
rect 5054 53286 5066 53338
rect 5066 53286 5096 53338
rect 5120 53286 5130 53338
rect 5130 53286 5176 53338
rect 4880 53284 4936 53286
rect 4960 53284 5016 53286
rect 5040 53284 5096 53286
rect 5120 53284 5176 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4880 52250 4936 52252
rect 4960 52250 5016 52252
rect 5040 52250 5096 52252
rect 5120 52250 5176 52252
rect 4880 52198 4926 52250
rect 4926 52198 4936 52250
rect 4960 52198 4990 52250
rect 4990 52198 5002 52250
rect 5002 52198 5016 52250
rect 5040 52198 5054 52250
rect 5054 52198 5066 52250
rect 5066 52198 5096 52250
rect 5120 52198 5130 52250
rect 5130 52198 5176 52250
rect 4880 52196 4936 52198
rect 4960 52196 5016 52198
rect 5040 52196 5096 52198
rect 5120 52196 5176 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4880 51162 4936 51164
rect 4960 51162 5016 51164
rect 5040 51162 5096 51164
rect 5120 51162 5176 51164
rect 4880 51110 4926 51162
rect 4926 51110 4936 51162
rect 4960 51110 4990 51162
rect 4990 51110 5002 51162
rect 5002 51110 5016 51162
rect 5040 51110 5054 51162
rect 5054 51110 5066 51162
rect 5066 51110 5096 51162
rect 5120 51110 5130 51162
rect 5130 51110 5176 51162
rect 4880 51108 4936 51110
rect 4960 51108 5016 51110
rect 5040 51108 5096 51110
rect 5120 51108 5176 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4880 50074 4936 50076
rect 4960 50074 5016 50076
rect 5040 50074 5096 50076
rect 5120 50074 5176 50076
rect 4880 50022 4926 50074
rect 4926 50022 4936 50074
rect 4960 50022 4990 50074
rect 4990 50022 5002 50074
rect 5002 50022 5016 50074
rect 5040 50022 5054 50074
rect 5054 50022 5066 50074
rect 5066 50022 5096 50074
rect 5120 50022 5130 50074
rect 5130 50022 5176 50074
rect 4880 50020 4936 50022
rect 4960 50020 5016 50022
rect 5040 50020 5096 50022
rect 5120 50020 5176 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4880 48986 4936 48988
rect 4960 48986 5016 48988
rect 5040 48986 5096 48988
rect 5120 48986 5176 48988
rect 4880 48934 4926 48986
rect 4926 48934 4936 48986
rect 4960 48934 4990 48986
rect 4990 48934 5002 48986
rect 5002 48934 5016 48986
rect 5040 48934 5054 48986
rect 5054 48934 5066 48986
rect 5066 48934 5096 48986
rect 5120 48934 5130 48986
rect 5130 48934 5176 48986
rect 4880 48932 4936 48934
rect 4960 48932 5016 48934
rect 5040 48932 5096 48934
rect 5120 48932 5176 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4880 47898 4936 47900
rect 4960 47898 5016 47900
rect 5040 47898 5096 47900
rect 5120 47898 5176 47900
rect 4880 47846 4926 47898
rect 4926 47846 4936 47898
rect 4960 47846 4990 47898
rect 4990 47846 5002 47898
rect 5002 47846 5016 47898
rect 5040 47846 5054 47898
rect 5054 47846 5066 47898
rect 5066 47846 5096 47898
rect 5120 47846 5130 47898
rect 5130 47846 5176 47898
rect 4880 47844 4936 47846
rect 4960 47844 5016 47846
rect 5040 47844 5096 47846
rect 5120 47844 5176 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4880 46810 4936 46812
rect 4960 46810 5016 46812
rect 5040 46810 5096 46812
rect 5120 46810 5176 46812
rect 4880 46758 4926 46810
rect 4926 46758 4936 46810
rect 4960 46758 4990 46810
rect 4990 46758 5002 46810
rect 5002 46758 5016 46810
rect 5040 46758 5054 46810
rect 5054 46758 5066 46810
rect 5066 46758 5096 46810
rect 5120 46758 5130 46810
rect 5130 46758 5176 46810
rect 4880 46756 4936 46758
rect 4960 46756 5016 46758
rect 5040 46756 5096 46758
rect 5120 46756 5176 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4880 45722 4936 45724
rect 4960 45722 5016 45724
rect 5040 45722 5096 45724
rect 5120 45722 5176 45724
rect 4880 45670 4926 45722
rect 4926 45670 4936 45722
rect 4960 45670 4990 45722
rect 4990 45670 5002 45722
rect 5002 45670 5016 45722
rect 5040 45670 5054 45722
rect 5054 45670 5066 45722
rect 5066 45670 5096 45722
rect 5120 45670 5130 45722
rect 5130 45670 5176 45722
rect 4880 45668 4936 45670
rect 4960 45668 5016 45670
rect 5040 45668 5096 45670
rect 5120 45668 5176 45670
rect 1674 30640 1730 30696
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4880 44634 4936 44636
rect 4960 44634 5016 44636
rect 5040 44634 5096 44636
rect 5120 44634 5176 44636
rect 4880 44582 4926 44634
rect 4926 44582 4936 44634
rect 4960 44582 4990 44634
rect 4990 44582 5002 44634
rect 5002 44582 5016 44634
rect 5040 44582 5054 44634
rect 5054 44582 5066 44634
rect 5066 44582 5096 44634
rect 5120 44582 5130 44634
rect 5130 44582 5176 44634
rect 4880 44580 4936 44582
rect 4960 44580 5016 44582
rect 5040 44580 5096 44582
rect 5120 44580 5176 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 35600 54426 35656 54428
rect 35680 54426 35736 54428
rect 35760 54426 35816 54428
rect 35840 54426 35896 54428
rect 35600 54374 35646 54426
rect 35646 54374 35656 54426
rect 35680 54374 35710 54426
rect 35710 54374 35722 54426
rect 35722 54374 35736 54426
rect 35760 54374 35774 54426
rect 35774 54374 35786 54426
rect 35786 54374 35816 54426
rect 35840 54374 35850 54426
rect 35850 54374 35896 54426
rect 35600 54372 35656 54374
rect 35680 54372 35736 54374
rect 35760 54372 35816 54374
rect 35840 54372 35896 54374
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 35600 53338 35656 53340
rect 35680 53338 35736 53340
rect 35760 53338 35816 53340
rect 35840 53338 35896 53340
rect 35600 53286 35646 53338
rect 35646 53286 35656 53338
rect 35680 53286 35710 53338
rect 35710 53286 35722 53338
rect 35722 53286 35736 53338
rect 35760 53286 35774 53338
rect 35774 53286 35786 53338
rect 35786 53286 35816 53338
rect 35840 53286 35850 53338
rect 35850 53286 35896 53338
rect 35600 53284 35656 53286
rect 35680 53284 35736 53286
rect 35760 53284 35816 53286
rect 35840 53284 35896 53286
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 35600 52250 35656 52252
rect 35680 52250 35736 52252
rect 35760 52250 35816 52252
rect 35840 52250 35896 52252
rect 35600 52198 35646 52250
rect 35646 52198 35656 52250
rect 35680 52198 35710 52250
rect 35710 52198 35722 52250
rect 35722 52198 35736 52250
rect 35760 52198 35774 52250
rect 35774 52198 35786 52250
rect 35786 52198 35816 52250
rect 35840 52198 35850 52250
rect 35850 52198 35896 52250
rect 35600 52196 35656 52198
rect 35680 52196 35736 52198
rect 35760 52196 35816 52198
rect 35840 52196 35896 52198
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 35600 51162 35656 51164
rect 35680 51162 35736 51164
rect 35760 51162 35816 51164
rect 35840 51162 35896 51164
rect 35600 51110 35646 51162
rect 35646 51110 35656 51162
rect 35680 51110 35710 51162
rect 35710 51110 35722 51162
rect 35722 51110 35736 51162
rect 35760 51110 35774 51162
rect 35774 51110 35786 51162
rect 35786 51110 35816 51162
rect 35840 51110 35850 51162
rect 35850 51110 35896 51162
rect 35600 51108 35656 51110
rect 35680 51108 35736 51110
rect 35760 51108 35816 51110
rect 35840 51108 35896 51110
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 35600 50074 35656 50076
rect 35680 50074 35736 50076
rect 35760 50074 35816 50076
rect 35840 50074 35896 50076
rect 35600 50022 35646 50074
rect 35646 50022 35656 50074
rect 35680 50022 35710 50074
rect 35710 50022 35722 50074
rect 35722 50022 35736 50074
rect 35760 50022 35774 50074
rect 35774 50022 35786 50074
rect 35786 50022 35816 50074
rect 35840 50022 35850 50074
rect 35850 50022 35896 50074
rect 35600 50020 35656 50022
rect 35680 50020 35736 50022
rect 35760 50020 35816 50022
rect 35840 50020 35896 50022
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 35600 48986 35656 48988
rect 35680 48986 35736 48988
rect 35760 48986 35816 48988
rect 35840 48986 35896 48988
rect 35600 48934 35646 48986
rect 35646 48934 35656 48986
rect 35680 48934 35710 48986
rect 35710 48934 35722 48986
rect 35722 48934 35736 48986
rect 35760 48934 35774 48986
rect 35774 48934 35786 48986
rect 35786 48934 35816 48986
rect 35840 48934 35850 48986
rect 35850 48934 35896 48986
rect 35600 48932 35656 48934
rect 35680 48932 35736 48934
rect 35760 48932 35816 48934
rect 35840 48932 35896 48934
rect 31206 38528 31262 38584
rect 32954 45736 33010 45792
rect 31850 40976 31906 41032
rect 31758 38528 31814 38584
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 35600 47898 35656 47900
rect 35680 47898 35736 47900
rect 35760 47898 35816 47900
rect 35840 47898 35896 47900
rect 35600 47846 35646 47898
rect 35646 47846 35656 47898
rect 35680 47846 35710 47898
rect 35710 47846 35722 47898
rect 35722 47846 35736 47898
rect 35760 47846 35774 47898
rect 35774 47846 35786 47898
rect 35786 47846 35816 47898
rect 35840 47846 35850 47898
rect 35850 47846 35896 47898
rect 35600 47844 35656 47846
rect 35680 47844 35736 47846
rect 35760 47844 35816 47846
rect 35840 47844 35896 47846
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 35600 46810 35656 46812
rect 35680 46810 35736 46812
rect 35760 46810 35816 46812
rect 35840 46810 35896 46812
rect 35600 46758 35646 46810
rect 35646 46758 35656 46810
rect 35680 46758 35710 46810
rect 35710 46758 35722 46810
rect 35722 46758 35736 46810
rect 35760 46758 35774 46810
rect 35774 46758 35786 46810
rect 35786 46758 35816 46810
rect 35840 46758 35850 46810
rect 35850 46758 35896 46810
rect 35600 46756 35656 46758
rect 35680 46756 35736 46758
rect 35760 46756 35816 46758
rect 35840 46756 35896 46758
rect 35600 45722 35656 45724
rect 35680 45722 35736 45724
rect 35760 45722 35816 45724
rect 35840 45722 35896 45724
rect 35600 45670 35646 45722
rect 35646 45670 35656 45722
rect 35680 45670 35710 45722
rect 35710 45670 35722 45722
rect 35722 45670 35736 45722
rect 35760 45670 35774 45722
rect 35774 45670 35786 45722
rect 35786 45670 35816 45722
rect 35840 45670 35850 45722
rect 35850 45670 35896 45722
rect 35600 45668 35656 45670
rect 35680 45668 35736 45670
rect 35760 45668 35816 45670
rect 35840 45668 35896 45670
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 32678 38528 32734 38584
rect 34150 41964 34152 41984
rect 34152 41964 34204 41984
rect 34204 41964 34206 41984
rect 34150 41928 34206 41964
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 33322 36100 33378 36136
rect 33322 36080 33324 36100
rect 33324 36080 33376 36100
rect 33376 36080 33378 36100
rect 33690 38800 33746 38856
rect 33690 36624 33746 36680
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 35600 44634 35656 44636
rect 35680 44634 35736 44636
rect 35760 44634 35816 44636
rect 35840 44634 35896 44636
rect 35600 44582 35646 44634
rect 35646 44582 35656 44634
rect 35680 44582 35710 44634
rect 35710 44582 35722 44634
rect 35722 44582 35736 44634
rect 35760 44582 35774 44634
rect 35774 44582 35786 44634
rect 35786 44582 35816 44634
rect 35840 44582 35850 44634
rect 35850 44582 35896 44634
rect 35600 44580 35656 44582
rect 35680 44580 35736 44582
rect 35760 44580 35816 44582
rect 35840 44580 35896 44582
rect 35600 43546 35656 43548
rect 35680 43546 35736 43548
rect 35760 43546 35816 43548
rect 35840 43546 35896 43548
rect 35600 43494 35646 43546
rect 35646 43494 35656 43546
rect 35680 43494 35710 43546
rect 35710 43494 35722 43546
rect 35722 43494 35736 43546
rect 35760 43494 35774 43546
rect 35774 43494 35786 43546
rect 35786 43494 35816 43546
rect 35840 43494 35850 43546
rect 35850 43494 35896 43546
rect 35600 43492 35656 43494
rect 35680 43492 35736 43494
rect 35760 43492 35816 43494
rect 35840 43492 35896 43494
rect 36082 43288 36138 43344
rect 35600 42458 35656 42460
rect 35680 42458 35736 42460
rect 35760 42458 35816 42460
rect 35840 42458 35896 42460
rect 35600 42406 35646 42458
rect 35646 42406 35656 42458
rect 35680 42406 35710 42458
rect 35710 42406 35722 42458
rect 35722 42406 35736 42458
rect 35760 42406 35774 42458
rect 35774 42406 35786 42458
rect 35786 42406 35816 42458
rect 35840 42406 35850 42458
rect 35850 42406 35896 42458
rect 35600 42404 35656 42406
rect 35680 42404 35736 42406
rect 35760 42404 35816 42406
rect 35840 42404 35896 42406
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 35600 41370 35656 41372
rect 35680 41370 35736 41372
rect 35760 41370 35816 41372
rect 35840 41370 35896 41372
rect 35600 41318 35646 41370
rect 35646 41318 35656 41370
rect 35680 41318 35710 41370
rect 35710 41318 35722 41370
rect 35722 41318 35736 41370
rect 35760 41318 35774 41370
rect 35774 41318 35786 41370
rect 35786 41318 35816 41370
rect 35840 41318 35850 41370
rect 35850 41318 35896 41370
rect 35600 41316 35656 41318
rect 35680 41316 35736 41318
rect 35760 41316 35816 41318
rect 35840 41316 35896 41318
rect 35806 40976 35862 41032
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 33782 35944 33838 36000
rect 35600 40282 35656 40284
rect 35680 40282 35736 40284
rect 35760 40282 35816 40284
rect 35840 40282 35896 40284
rect 35600 40230 35646 40282
rect 35646 40230 35656 40282
rect 35680 40230 35710 40282
rect 35710 40230 35722 40282
rect 35722 40230 35736 40282
rect 35760 40230 35774 40282
rect 35774 40230 35786 40282
rect 35786 40230 35816 40282
rect 35840 40230 35850 40282
rect 35850 40230 35896 40282
rect 35600 40228 35656 40230
rect 35680 40228 35736 40230
rect 35760 40228 35816 40230
rect 35840 40228 35896 40230
rect 35600 39194 35656 39196
rect 35680 39194 35736 39196
rect 35760 39194 35816 39196
rect 35840 39194 35896 39196
rect 35600 39142 35646 39194
rect 35646 39142 35656 39194
rect 35680 39142 35710 39194
rect 35710 39142 35722 39194
rect 35722 39142 35736 39194
rect 35760 39142 35774 39194
rect 35774 39142 35786 39194
rect 35786 39142 35816 39194
rect 35840 39142 35850 39194
rect 35850 39142 35896 39194
rect 35600 39140 35656 39142
rect 35680 39140 35736 39142
rect 35760 39140 35816 39142
rect 35840 39140 35896 39142
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 35600 38106 35656 38108
rect 35680 38106 35736 38108
rect 35760 38106 35816 38108
rect 35840 38106 35896 38108
rect 35600 38054 35646 38106
rect 35646 38054 35656 38106
rect 35680 38054 35710 38106
rect 35710 38054 35722 38106
rect 35722 38054 35736 38106
rect 35760 38054 35774 38106
rect 35774 38054 35786 38106
rect 35786 38054 35816 38106
rect 35840 38054 35850 38106
rect 35850 38054 35896 38106
rect 35600 38052 35656 38054
rect 35680 38052 35736 38054
rect 35760 38052 35816 38054
rect 35840 38052 35896 38054
rect 31298 29144 31354 29200
rect 32402 30232 32458 30288
rect 34334 30776 34390 30832
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 35898 36624 35954 36680
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 34334 28192 34390 28248
rect 35346 30368 35402 30424
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 35346 29688 35402 29744
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 36726 43308 36782 43344
rect 36726 43288 36728 43308
rect 36728 43288 36780 43308
rect 36780 43288 36782 43308
rect 36542 38256 36598 38312
rect 36634 36080 36690 36136
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 36358 29180 36360 29200
rect 36360 29180 36412 29200
rect 36412 29180 36414 29200
rect 36358 29144 36414 29180
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 38014 44784 38070 44840
rect 37554 40704 37610 40760
rect 37738 40160 37794 40216
rect 37646 39888 37702 39944
rect 38106 40180 38162 40216
rect 38106 40160 38108 40180
rect 38108 40160 38160 40180
rect 38160 40160 38162 40180
rect 38106 39924 38108 39944
rect 38108 39924 38160 39944
rect 38160 39924 38162 39944
rect 38106 39888 38162 39924
rect 38106 38800 38162 38856
rect 38106 38292 38108 38312
rect 38108 38292 38160 38312
rect 38160 38292 38162 38312
rect 38106 38256 38162 38292
rect 38106 36624 38162 36680
rect 38566 41268 38622 41304
rect 38566 41248 38568 41268
rect 38568 41248 38620 41268
rect 38620 41248 38622 41268
rect 38382 41132 38438 41168
rect 39210 43308 39266 43344
rect 39210 43288 39212 43308
rect 39212 43288 39264 43308
rect 39264 43288 39266 43308
rect 40498 45484 40554 45520
rect 40498 45464 40500 45484
rect 40500 45464 40552 45484
rect 40552 45464 40554 45484
rect 40406 43696 40462 43752
rect 40314 43308 40370 43344
rect 40314 43288 40316 43308
rect 40316 43288 40368 43308
rect 40368 43288 40370 43308
rect 38382 41112 38384 41132
rect 38384 41112 38436 41132
rect 38436 41112 38438 41132
rect 38566 40996 38622 41032
rect 38566 40976 38568 40996
rect 38568 40976 38620 40996
rect 38620 40976 38622 40996
rect 37278 32544 37334 32600
rect 37554 32564 37610 32600
rect 37554 32544 37556 32564
rect 37556 32544 37608 32564
rect 37608 32544 37610 32564
rect 37094 29416 37150 29472
rect 37830 32000 37886 32056
rect 39302 34720 39358 34776
rect 38382 32544 38438 32600
rect 38658 32428 38714 32464
rect 38658 32408 38660 32428
rect 38660 32408 38712 32428
rect 38712 32408 38714 32428
rect 38382 32272 38438 32328
rect 38198 29996 38200 30016
rect 38200 29996 38252 30016
rect 38252 29996 38254 30016
rect 38198 29960 38254 29996
rect 38658 32136 38714 32192
rect 38566 32020 38622 32056
rect 38566 32000 38568 32020
rect 38568 32000 38620 32020
rect 38620 32000 38622 32020
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 40222 41556 40224 41576
rect 40224 41556 40276 41576
rect 40276 41556 40278 41576
rect 40222 41520 40278 41556
rect 39946 39516 39948 39536
rect 39948 39516 40000 39536
rect 40000 39516 40002 39536
rect 39946 39480 40002 39516
rect 39026 30132 39028 30152
rect 39028 30132 39080 30152
rect 39080 30132 39082 30152
rect 39026 30096 39082 30132
rect 39210 29300 39266 29336
rect 39210 29280 39212 29300
rect 39212 29280 39264 29300
rect 39264 29280 39266 29300
rect 39486 28056 39542 28112
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 39026 24148 39028 24168
rect 39028 24148 39080 24168
rect 39080 24148 39082 24168
rect 39026 24112 39082 24148
rect 40406 29824 40462 29880
rect 40498 29008 40554 29064
rect 40314 28872 40370 28928
rect 41050 43172 41106 43208
rect 41050 43152 41052 43172
rect 41052 43152 41104 43172
rect 41104 43152 41106 43172
rect 41142 43016 41198 43072
rect 40958 42880 41014 42936
rect 41878 47404 41880 47424
rect 41880 47404 41932 47424
rect 41932 47404 41934 47424
rect 41878 47368 41934 47404
rect 41510 43052 41512 43072
rect 41512 43052 41564 43072
rect 41564 43052 41566 43072
rect 41510 43016 41566 43052
rect 42154 43152 42210 43208
rect 41326 41556 41328 41576
rect 41328 41556 41380 41576
rect 41380 41556 41382 41576
rect 41326 41520 41382 41556
rect 42154 39516 42156 39536
rect 42156 39516 42208 39536
rect 42208 39516 42210 39536
rect 42154 39480 42210 39516
rect 41878 33108 41934 33144
rect 41878 33088 41880 33108
rect 41880 33088 41932 33108
rect 41932 33088 41934 33108
rect 41326 30368 41382 30424
rect 41050 29688 41106 29744
rect 41050 29552 41106 29608
rect 40682 28328 40738 28384
rect 40958 29144 41014 29200
rect 41142 29300 41198 29336
rect 41142 29280 41144 29300
rect 41144 29280 41196 29300
rect 41196 29280 41198 29300
rect 41602 30096 41658 30152
rect 41510 29824 41566 29880
rect 41234 28872 41290 28928
rect 40130 26560 40186 26616
rect 41234 28328 41290 28384
rect 41418 28328 41474 28384
rect 42798 37984 42854 38040
rect 44638 45464 44694 45520
rect 45374 43732 45376 43752
rect 45376 43732 45428 43752
rect 45428 43732 45430 43752
rect 45374 43696 45430 43732
rect 42522 28076 42578 28112
rect 42522 28056 42524 28076
rect 42524 28056 42576 28076
rect 42576 28056 42578 28076
rect 43810 34720 43866 34776
rect 42706 31204 42762 31240
rect 42706 31184 42708 31204
rect 42708 31184 42760 31204
rect 42760 31184 42762 31204
rect 42706 29688 42762 29744
rect 42982 29960 43038 30016
rect 41602 24148 41604 24168
rect 41604 24148 41656 24168
rect 41656 24148 41658 24168
rect 41602 24112 41658 24148
rect 43994 29588 43996 29608
rect 43996 29588 44048 29608
rect 44048 29588 44050 29608
rect 43994 29552 44050 29588
rect 44270 29144 44326 29200
rect 46202 45892 46258 45928
rect 46202 45872 46204 45892
rect 46204 45872 46256 45892
rect 46256 45872 46258 45892
rect 48778 45600 48834 45656
rect 48318 39924 48320 39944
rect 48320 39924 48372 39944
rect 48372 39924 48374 39944
rect 48318 39888 48374 39924
rect 45926 31864 45982 31920
rect 45374 31320 45430 31376
rect 45098 29416 45154 29472
rect 45466 29416 45522 29472
rect 45558 27240 45614 27296
rect 45834 29280 45890 29336
rect 45926 28872 45982 28928
rect 47398 33088 47454 33144
rect 46754 30676 46756 30696
rect 46756 30676 46808 30696
rect 46808 30676 46810 30696
rect 46754 30640 46810 30676
rect 46938 31340 46994 31376
rect 46938 31320 46940 31340
rect 46940 31320 46992 31340
rect 46992 31320 46994 31340
rect 46846 30368 46902 30424
rect 47030 30776 47086 30832
rect 47214 29416 47270 29472
rect 47122 28872 47178 28928
rect 47582 30368 47638 30424
rect 46662 26560 46718 26616
rect 46938 26036 46994 26072
rect 46938 26016 46940 26036
rect 46940 26016 46992 26036
rect 46992 26016 46994 26036
rect 48226 37984 48282 38040
rect 49330 42628 49386 42664
rect 49330 42608 49332 42628
rect 49332 42608 49384 42628
rect 49384 42608 49386 42628
rect 49238 42508 49240 42528
rect 49240 42508 49292 42528
rect 49292 42508 49294 42528
rect 49238 42472 49294 42508
rect 49146 41384 49202 41440
rect 49606 41384 49662 41440
rect 49330 37984 49386 38040
rect 50342 42628 50398 42664
rect 50342 42608 50344 42628
rect 50344 42608 50396 42628
rect 50396 42608 50398 42628
rect 49974 38392 50030 38448
rect 47858 29280 47914 29336
rect 47950 29164 48006 29200
rect 47950 29144 47952 29164
rect 47952 29144 48004 29164
rect 48004 29144 48006 29164
rect 48134 30660 48190 30696
rect 48134 30640 48136 30660
rect 48136 30640 48188 30660
rect 48188 30640 48190 30660
rect 48226 29144 48282 29200
rect 47950 27648 48006 27704
rect 48962 28076 49018 28112
rect 48962 28056 48964 28076
rect 48964 28056 49016 28076
rect 49016 28056 49018 28076
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 49606 28212 49662 28248
rect 49606 28192 49608 28212
rect 49608 28192 49660 28212
rect 49660 28192 49662 28212
rect 51998 42472 52054 42528
rect 50802 38392 50858 38448
rect 50342 29144 50398 29200
rect 52826 38392 52882 38448
rect 51998 28212 52054 28248
rect 51998 28192 52000 28212
rect 52000 28192 52052 28212
rect 52052 28192 52054 28212
rect 51078 28056 51134 28112
rect 51906 27648 51962 27704
rect 51630 27512 51686 27568
rect 53102 27668 53158 27704
rect 53102 27648 53104 27668
rect 53104 27648 53156 27668
rect 53156 27648 53158 27668
rect 53378 29144 53434 29200
rect 55402 29164 55458 29200
rect 55402 29144 55404 29164
rect 55404 29144 55456 29164
rect 55456 29144 55458 29164
rect 58254 29280 58310 29336
rect 58622 31184 58678 31240
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
<< metal3 >>
rect 4870 57696 5186 57697
rect 4870 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5186 57696
rect 4870 57631 5186 57632
rect 35590 57696 35906 57697
rect 35590 57632 35596 57696
rect 35660 57632 35676 57696
rect 35740 57632 35756 57696
rect 35820 57632 35836 57696
rect 35900 57632 35906 57696
rect 35590 57631 35906 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 4870 56608 5186 56609
rect 4870 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5186 56608
rect 4870 56543 5186 56544
rect 35590 56608 35906 56609
rect 35590 56544 35596 56608
rect 35660 56544 35676 56608
rect 35740 56544 35756 56608
rect 35820 56544 35836 56608
rect 35900 56544 35906 56608
rect 35590 56543 35906 56544
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 4870 55520 5186 55521
rect 4870 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5186 55520
rect 4870 55455 5186 55456
rect 35590 55520 35906 55521
rect 35590 55456 35596 55520
rect 35660 55456 35676 55520
rect 35740 55456 35756 55520
rect 35820 55456 35836 55520
rect 35900 55456 35906 55520
rect 35590 55455 35906 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 4870 54432 5186 54433
rect 4870 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5186 54432
rect 4870 54367 5186 54368
rect 35590 54432 35906 54433
rect 35590 54368 35596 54432
rect 35660 54368 35676 54432
rect 35740 54368 35756 54432
rect 35820 54368 35836 54432
rect 35900 54368 35906 54432
rect 35590 54367 35906 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 4870 53344 5186 53345
rect 4870 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5186 53344
rect 4870 53279 5186 53280
rect 35590 53344 35906 53345
rect 35590 53280 35596 53344
rect 35660 53280 35676 53344
rect 35740 53280 35756 53344
rect 35820 53280 35836 53344
rect 35900 53280 35906 53344
rect 35590 53279 35906 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 4870 52256 5186 52257
rect 4870 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5186 52256
rect 4870 52191 5186 52192
rect 35590 52256 35906 52257
rect 35590 52192 35596 52256
rect 35660 52192 35676 52256
rect 35740 52192 35756 52256
rect 35820 52192 35836 52256
rect 35900 52192 35906 52256
rect 35590 52191 35906 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 4870 51168 5186 51169
rect 4870 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5186 51168
rect 4870 51103 5186 51104
rect 35590 51168 35906 51169
rect 35590 51104 35596 51168
rect 35660 51104 35676 51168
rect 35740 51104 35756 51168
rect 35820 51104 35836 51168
rect 35900 51104 35906 51168
rect 35590 51103 35906 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 4870 50080 5186 50081
rect 4870 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5186 50080
rect 4870 50015 5186 50016
rect 35590 50080 35906 50081
rect 35590 50016 35596 50080
rect 35660 50016 35676 50080
rect 35740 50016 35756 50080
rect 35820 50016 35836 50080
rect 35900 50016 35906 50080
rect 35590 50015 35906 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 4870 48992 5186 48993
rect 4870 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5186 48992
rect 4870 48927 5186 48928
rect 35590 48992 35906 48993
rect 35590 48928 35596 48992
rect 35660 48928 35676 48992
rect 35740 48928 35756 48992
rect 35820 48928 35836 48992
rect 35900 48928 35906 48992
rect 35590 48927 35906 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 4870 47904 5186 47905
rect 4870 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5186 47904
rect 4870 47839 5186 47840
rect 35590 47904 35906 47905
rect 35590 47840 35596 47904
rect 35660 47840 35676 47904
rect 35740 47840 35756 47904
rect 35820 47840 35836 47904
rect 35900 47840 35906 47904
rect 35590 47839 35906 47840
rect 41873 47426 41939 47429
rect 42006 47426 42012 47428
rect 41873 47424 42012 47426
rect 41873 47368 41878 47424
rect 41934 47368 42012 47424
rect 41873 47366 42012 47368
rect 41873 47363 41939 47366
rect 42006 47364 42012 47366
rect 42076 47364 42082 47428
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 4870 46816 5186 46817
rect 4870 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5186 46816
rect 4870 46751 5186 46752
rect 35590 46816 35906 46817
rect 35590 46752 35596 46816
rect 35660 46752 35676 46816
rect 35740 46752 35756 46816
rect 35820 46752 35836 46816
rect 35900 46752 35906 46816
rect 35590 46751 35906 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 42006 45868 42012 45932
rect 42076 45930 42082 45932
rect 46197 45930 46263 45933
rect 42076 45928 46263 45930
rect 42076 45872 46202 45928
rect 46258 45872 46263 45928
rect 42076 45870 46263 45872
rect 42076 45868 42082 45870
rect 46197 45867 46263 45870
rect 32438 45732 32444 45796
rect 32508 45794 32514 45796
rect 32949 45794 33015 45797
rect 32508 45792 33015 45794
rect 32508 45736 32954 45792
rect 33010 45736 33015 45792
rect 32508 45734 33015 45736
rect 32508 45732 32514 45734
rect 32949 45731 33015 45734
rect 4870 45728 5186 45729
rect 4870 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5186 45728
rect 4870 45663 5186 45664
rect 35590 45728 35906 45729
rect 35590 45664 35596 45728
rect 35660 45664 35676 45728
rect 35740 45664 35756 45728
rect 35820 45664 35836 45728
rect 35900 45664 35906 45728
rect 35590 45663 35906 45664
rect 48630 45596 48636 45660
rect 48700 45658 48706 45660
rect 48773 45658 48839 45661
rect 48700 45656 48839 45658
rect 48700 45600 48778 45656
rect 48834 45600 48839 45656
rect 48700 45598 48839 45600
rect 48700 45596 48706 45598
rect 48773 45595 48839 45598
rect 40493 45522 40559 45525
rect 44633 45522 44699 45525
rect 40493 45520 44699 45522
rect 40493 45464 40498 45520
rect 40554 45464 44638 45520
rect 44694 45464 44699 45520
rect 40493 45462 44699 45464
rect 40493 45459 40559 45462
rect 44633 45459 44699 45462
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 37590 44780 37596 44844
rect 37660 44842 37666 44844
rect 38009 44842 38075 44845
rect 37660 44840 38075 44842
rect 37660 44784 38014 44840
rect 38070 44784 38075 44840
rect 37660 44782 38075 44784
rect 37660 44780 37666 44782
rect 38009 44779 38075 44782
rect 4870 44640 5186 44641
rect 4870 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5186 44640
rect 4870 44575 5186 44576
rect 35590 44640 35906 44641
rect 35590 44576 35596 44640
rect 35660 44576 35676 44640
rect 35740 44576 35756 44640
rect 35820 44576 35836 44640
rect 35900 44576 35906 44640
rect 35590 44575 35906 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 40401 43754 40467 43757
rect 45369 43754 45435 43757
rect 40401 43752 45435 43754
rect 40401 43696 40406 43752
rect 40462 43696 45374 43752
rect 45430 43696 45435 43752
rect 40401 43694 45435 43696
rect 40401 43691 40467 43694
rect 45369 43691 45435 43694
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 35590 43552 35906 43553
rect 35590 43488 35596 43552
rect 35660 43488 35676 43552
rect 35740 43488 35756 43552
rect 35820 43488 35836 43552
rect 35900 43488 35906 43552
rect 35590 43487 35906 43488
rect 36077 43346 36143 43349
rect 36721 43346 36787 43349
rect 36077 43344 36787 43346
rect 36077 43288 36082 43344
rect 36138 43288 36726 43344
rect 36782 43288 36787 43344
rect 36077 43286 36787 43288
rect 36077 43283 36143 43286
rect 36721 43283 36787 43286
rect 39205 43346 39271 43349
rect 40309 43346 40375 43349
rect 39205 43344 40375 43346
rect 39205 43288 39210 43344
rect 39266 43288 40314 43344
rect 40370 43288 40375 43344
rect 39205 43286 40375 43288
rect 39205 43283 39271 43286
rect 40309 43283 40375 43286
rect 41045 43210 41111 43213
rect 42149 43210 42215 43213
rect 41045 43208 42215 43210
rect 41045 43152 41050 43208
rect 41106 43152 42154 43208
rect 42210 43152 42215 43208
rect 41045 43150 42215 43152
rect 41045 43147 41111 43150
rect 42149 43147 42215 43150
rect 41137 43074 41203 43077
rect 41505 43074 41571 43077
rect 41137 43072 41571 43074
rect 41137 43016 41142 43072
rect 41198 43016 41510 43072
rect 41566 43016 41571 43072
rect 41137 43014 41571 43016
rect 41137 43011 41203 43014
rect 41505 43011 41571 43014
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 40953 42938 41019 42941
rect 41086 42938 41092 42940
rect 40953 42936 41092 42938
rect 40953 42880 40958 42936
rect 41014 42880 41092 42936
rect 40953 42878 41092 42880
rect 40953 42875 41019 42878
rect 41086 42876 41092 42878
rect 41156 42876 41162 42940
rect 49325 42666 49391 42669
rect 50337 42666 50403 42669
rect 49325 42664 50403 42666
rect 49325 42608 49330 42664
rect 49386 42608 50342 42664
rect 50398 42608 50403 42664
rect 49325 42606 50403 42608
rect 49325 42603 49391 42606
rect 50337 42603 50403 42606
rect 49233 42530 49299 42533
rect 51993 42530 52059 42533
rect 49233 42528 52059 42530
rect 49233 42472 49238 42528
rect 49294 42472 51998 42528
rect 52054 42472 52059 42528
rect 49233 42470 52059 42472
rect 49233 42467 49299 42470
rect 51993 42467 52059 42470
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 35590 42464 35906 42465
rect 35590 42400 35596 42464
rect 35660 42400 35676 42464
rect 35740 42400 35756 42464
rect 35820 42400 35836 42464
rect 35900 42400 35906 42464
rect 35590 42399 35906 42400
rect 34145 41986 34211 41989
rect 34278 41986 34284 41988
rect 34145 41984 34284 41986
rect 34145 41928 34150 41984
rect 34206 41928 34284 41984
rect 34145 41926 34284 41928
rect 34145 41923 34211 41926
rect 34278 41924 34284 41926
rect 34348 41924 34354 41988
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 40217 41578 40283 41581
rect 41321 41578 41387 41581
rect 40217 41576 41387 41578
rect 40217 41520 40222 41576
rect 40278 41520 41326 41576
rect 41382 41520 41387 41576
rect 40217 41518 41387 41520
rect 40217 41515 40283 41518
rect 41321 41515 41387 41518
rect 49141 41442 49207 41445
rect 49601 41442 49667 41445
rect 49141 41440 49667 41442
rect 49141 41384 49146 41440
rect 49202 41384 49606 41440
rect 49662 41384 49667 41440
rect 49141 41382 49667 41384
rect 49141 41379 49207 41382
rect 49601 41379 49667 41382
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 35590 41376 35906 41377
rect 35590 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35906 41376
rect 35590 41311 35906 41312
rect 38561 41308 38627 41309
rect 38510 41306 38516 41308
rect 38470 41246 38516 41306
rect 38580 41304 38627 41308
rect 38622 41248 38627 41304
rect 38510 41244 38516 41246
rect 38580 41244 38627 41248
rect 38518 41243 38627 41244
rect 38377 41170 38443 41173
rect 38518 41170 38578 41243
rect 38377 41168 38578 41170
rect 38377 41112 38382 41168
rect 38438 41112 38578 41168
rect 38377 41110 38578 41112
rect 38377 41107 38443 41110
rect 31845 41034 31911 41037
rect 35801 41034 35867 41037
rect 38561 41034 38627 41037
rect 31845 41032 38627 41034
rect 31845 40976 31850 41032
rect 31906 40976 35806 41032
rect 35862 40976 38566 41032
rect 38622 40976 38627 41032
rect 31845 40974 38627 40976
rect 31845 40971 31911 40974
rect 35801 40971 35867 40974
rect 38561 40971 38627 40974
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 37549 40762 37615 40765
rect 38510 40762 38516 40764
rect 37549 40760 38516 40762
rect 37549 40704 37554 40760
rect 37610 40704 38516 40760
rect 37549 40702 38516 40704
rect 37549 40699 37615 40702
rect 38510 40700 38516 40702
rect 38580 40700 38586 40764
rect 4870 40288 5186 40289
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 35590 40288 35906 40289
rect 35590 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35906 40288
rect 35590 40223 35906 40224
rect 37733 40218 37799 40221
rect 38101 40218 38167 40221
rect 37733 40216 38167 40218
rect 37733 40160 37738 40216
rect 37794 40160 38106 40216
rect 38162 40160 38167 40216
rect 37733 40158 38167 40160
rect 37733 40155 37799 40158
rect 38101 40155 38167 40158
rect 37641 39946 37707 39949
rect 38101 39946 38167 39949
rect 48313 39948 48379 39949
rect 37641 39944 38167 39946
rect 37641 39888 37646 39944
rect 37702 39888 38106 39944
rect 38162 39888 38167 39944
rect 37641 39886 38167 39888
rect 37641 39883 37707 39886
rect 38101 39883 38167 39886
rect 48262 39884 48268 39948
rect 48332 39946 48379 39948
rect 48630 39946 48636 39948
rect 48332 39944 48636 39946
rect 48374 39888 48636 39944
rect 48332 39886 48636 39888
rect 48332 39884 48379 39886
rect 48630 39884 48636 39886
rect 48700 39884 48706 39948
rect 48313 39883 48379 39884
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 39941 39538 40007 39541
rect 42149 39538 42215 39541
rect 39941 39536 42215 39538
rect 39941 39480 39946 39536
rect 40002 39480 42154 39536
rect 42210 39480 42215 39536
rect 39941 39478 42215 39480
rect 39941 39475 40007 39478
rect 42149 39475 42215 39478
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 35590 39200 35906 39201
rect 35590 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35906 39200
rect 35590 39135 35906 39136
rect 33685 38858 33751 38861
rect 38101 38858 38167 38861
rect 33685 38856 38167 38858
rect 33685 38800 33690 38856
rect 33746 38800 38106 38856
rect 38162 38800 38167 38856
rect 33685 38798 38167 38800
rect 33685 38795 33751 38798
rect 38101 38795 38167 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 31201 38586 31267 38589
rect 31753 38586 31819 38589
rect 32673 38586 32739 38589
rect 31201 38584 32739 38586
rect 31201 38528 31206 38584
rect 31262 38528 31758 38584
rect 31814 38528 32678 38584
rect 32734 38528 32739 38584
rect 31201 38526 32739 38528
rect 31201 38523 31267 38526
rect 31753 38523 31819 38526
rect 32673 38523 32739 38526
rect 49969 38450 50035 38453
rect 50797 38450 50863 38453
rect 52821 38450 52887 38453
rect 49969 38448 52887 38450
rect 49969 38392 49974 38448
rect 50030 38392 50802 38448
rect 50858 38392 52826 38448
rect 52882 38392 52887 38448
rect 49969 38390 52887 38392
rect 49969 38387 50035 38390
rect 50797 38387 50863 38390
rect 52821 38387 52887 38390
rect 36537 38314 36603 38317
rect 38101 38314 38167 38317
rect 36537 38312 38167 38314
rect 36537 38256 36542 38312
rect 36598 38256 38106 38312
rect 38162 38256 38167 38312
rect 36537 38254 38167 38256
rect 36537 38251 36603 38254
rect 38101 38251 38167 38254
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 35590 38112 35906 38113
rect 35590 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35906 38112
rect 35590 38047 35906 38048
rect 42793 38042 42859 38045
rect 48221 38042 48287 38045
rect 49325 38042 49391 38045
rect 42793 38040 49391 38042
rect 42793 37984 42798 38040
rect 42854 37984 48226 38040
rect 48282 37984 49330 38040
rect 49386 37984 49391 38040
rect 42793 37982 49391 37984
rect 42793 37979 42859 37982
rect 48221 37979 48287 37982
rect 49325 37979 49391 37982
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 33685 36682 33751 36685
rect 35893 36682 35959 36685
rect 38101 36682 38167 36685
rect 33685 36680 38167 36682
rect 33685 36624 33690 36680
rect 33746 36624 35898 36680
rect 35954 36624 38106 36680
rect 38162 36624 38167 36680
rect 33685 36622 38167 36624
rect 33685 36619 33751 36622
rect 35893 36619 35959 36622
rect 38101 36619 38167 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 33317 36138 33383 36141
rect 36629 36138 36695 36141
rect 33317 36136 36695 36138
rect 33317 36080 33322 36136
rect 33378 36080 36634 36136
rect 36690 36080 36695 36136
rect 33317 36078 36695 36080
rect 33317 36075 33383 36078
rect 33734 36005 33794 36078
rect 36629 36075 36695 36078
rect 33734 36000 33843 36005
rect 33734 35944 33782 36000
rect 33838 35944 33843 36000
rect 33734 35942 33843 35944
rect 33777 35939 33843 35942
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 39297 34778 39363 34781
rect 43805 34778 43871 34781
rect 39297 34776 43871 34778
rect 39297 34720 39302 34776
rect 39358 34720 43810 34776
rect 43866 34720 43871 34776
rect 39297 34718 43871 34720
rect 39297 34715 39363 34718
rect 43805 34715 43871 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 41873 33146 41939 33149
rect 42006 33146 42012 33148
rect 41873 33144 42012 33146
rect 41873 33088 41878 33144
rect 41934 33088 42012 33144
rect 41873 33086 42012 33088
rect 41873 33083 41939 33086
rect 42006 33084 42012 33086
rect 42076 33084 42082 33148
rect 47393 33146 47459 33149
rect 48262 33146 48268 33148
rect 47393 33144 48268 33146
rect 47393 33088 47398 33144
rect 47454 33088 48268 33144
rect 47393 33086 48268 33088
rect 47393 33083 47459 33086
rect 48262 33084 48268 33086
rect 48332 33084 48338 33148
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 37273 32602 37339 32605
rect 37549 32604 37615 32605
rect 37549 32602 37596 32604
rect 37273 32600 37596 32602
rect 37273 32544 37278 32600
rect 37334 32544 37554 32600
rect 37273 32542 37596 32544
rect 37273 32539 37339 32542
rect 37549 32540 37596 32542
rect 37660 32540 37666 32604
rect 38377 32602 38443 32605
rect 38334 32600 38443 32602
rect 38334 32544 38382 32600
rect 38438 32544 38443 32600
rect 37549 32539 37615 32540
rect 38334 32539 38443 32544
rect 38334 32333 38394 32539
rect 38653 32466 38719 32469
rect 38518 32464 38719 32466
rect 38518 32408 38658 32464
rect 38714 32408 38719 32464
rect 38518 32406 38719 32408
rect 38334 32328 38443 32333
rect 38334 32272 38382 32328
rect 38438 32272 38443 32328
rect 38334 32270 38443 32272
rect 38377 32267 38443 32270
rect 38518 32194 38578 32406
rect 38653 32403 38719 32406
rect 38653 32194 38719 32197
rect 38518 32192 38719 32194
rect 38518 32136 38658 32192
rect 38714 32136 38719 32192
rect 38518 32134 38719 32136
rect 38653 32131 38719 32134
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 37825 32058 37891 32061
rect 38561 32058 38627 32061
rect 37825 32056 38627 32058
rect 37825 32000 37830 32056
rect 37886 32000 38566 32056
rect 38622 32000 38627 32056
rect 37825 31998 38627 32000
rect 37825 31995 37891 31998
rect 38561 31995 38627 31998
rect 41086 31860 41092 31924
rect 41156 31922 41162 31924
rect 45921 31922 45987 31925
rect 41156 31920 45987 31922
rect 41156 31864 45926 31920
rect 45982 31864 45987 31920
rect 41156 31862 45987 31864
rect 41156 31860 41162 31862
rect 45921 31859 45987 31862
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 45369 31378 45435 31381
rect 46933 31378 46999 31381
rect 45369 31376 46999 31378
rect 45369 31320 45374 31376
rect 45430 31320 46938 31376
rect 46994 31320 46999 31376
rect 45369 31318 46999 31320
rect 45369 31315 45435 31318
rect 46933 31315 46999 31318
rect 42701 31242 42767 31245
rect 58617 31242 58683 31245
rect 42701 31240 58683 31242
rect 42701 31184 42706 31240
rect 42762 31184 58622 31240
rect 58678 31184 58683 31240
rect 42701 31182 58683 31184
rect 42701 31179 42767 31182
rect 58617 31179 58683 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 34329 30834 34395 30837
rect 47025 30834 47091 30837
rect 34329 30832 47091 30834
rect 34329 30776 34334 30832
rect 34390 30776 47030 30832
rect 47086 30776 47091 30832
rect 34329 30774 47091 30776
rect 34329 30771 34395 30774
rect 47025 30771 47091 30774
rect 200 30698 800 30728
rect 1669 30698 1735 30701
rect 200 30696 1735 30698
rect 200 30640 1674 30696
rect 1730 30640 1735 30696
rect 200 30638 1735 30640
rect 200 30608 800 30638
rect 1669 30635 1735 30638
rect 46749 30698 46815 30701
rect 48129 30698 48195 30701
rect 46749 30696 48195 30698
rect 46749 30640 46754 30696
rect 46810 30640 48134 30696
rect 48190 30640 48195 30696
rect 46749 30638 48195 30640
rect 46749 30635 46815 30638
rect 48129 30635 48195 30638
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 35341 30424 35407 30429
rect 35341 30368 35346 30424
rect 35402 30368 35407 30424
rect 35341 30363 35407 30368
rect 41321 30426 41387 30429
rect 46841 30426 46907 30429
rect 41321 30424 46907 30426
rect 41321 30368 41326 30424
rect 41382 30368 46846 30424
rect 46902 30368 46907 30424
rect 41321 30366 46907 30368
rect 41321 30363 41387 30366
rect 46841 30363 46907 30366
rect 47577 30426 47643 30429
rect 48262 30426 48268 30428
rect 47577 30424 48268 30426
rect 47577 30368 47582 30424
rect 47638 30368 48268 30424
rect 47577 30366 48268 30368
rect 47577 30363 47643 30366
rect 48262 30364 48268 30366
rect 48332 30364 48338 30428
rect 32397 30292 32463 30293
rect 32397 30290 32444 30292
rect 32352 30288 32444 30290
rect 32352 30232 32402 30288
rect 32352 30230 32444 30232
rect 32397 30228 32444 30230
rect 32508 30228 32514 30292
rect 32397 30227 32463 30228
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 35344 29749 35404 30363
rect 39021 30154 39087 30157
rect 41597 30154 41663 30157
rect 39021 30152 41663 30154
rect 39021 30096 39026 30152
rect 39082 30096 41602 30152
rect 41658 30096 41663 30152
rect 39021 30094 41663 30096
rect 39021 30091 39087 30094
rect 41597 30091 41663 30094
rect 38193 30018 38259 30021
rect 42977 30018 43043 30021
rect 38193 30016 43043 30018
rect 38193 29960 38198 30016
rect 38254 29960 42982 30016
rect 43038 29960 43043 30016
rect 38193 29958 43043 29960
rect 38193 29955 38259 29958
rect 42977 29955 43043 29958
rect 40401 29882 40467 29885
rect 41505 29882 41571 29885
rect 40401 29880 41571 29882
rect 40401 29824 40406 29880
rect 40462 29824 41510 29880
rect 41566 29824 41571 29880
rect 40401 29822 41571 29824
rect 40401 29819 40467 29822
rect 41505 29819 41571 29822
rect 35341 29744 35407 29749
rect 35341 29688 35346 29744
rect 35402 29688 35407 29744
rect 35341 29683 35407 29688
rect 41045 29746 41111 29749
rect 42701 29746 42767 29749
rect 41045 29744 42767 29746
rect 41045 29688 41050 29744
rect 41106 29688 42706 29744
rect 42762 29688 42767 29744
rect 41045 29686 42767 29688
rect 41045 29683 41111 29686
rect 42701 29683 42767 29686
rect 41045 29610 41111 29613
rect 43989 29610 44055 29613
rect 41045 29608 44055 29610
rect 41045 29552 41050 29608
rect 41106 29552 43994 29608
rect 44050 29552 44055 29608
rect 41045 29550 44055 29552
rect 41045 29547 41111 29550
rect 43989 29547 44055 29550
rect 37089 29474 37155 29477
rect 45093 29474 45159 29477
rect 37089 29472 45159 29474
rect 37089 29416 37094 29472
rect 37150 29416 45098 29472
rect 45154 29416 45159 29472
rect 37089 29414 45159 29416
rect 37089 29411 37155 29414
rect 45093 29411 45159 29414
rect 45461 29474 45527 29477
rect 46974 29474 46980 29476
rect 45461 29472 46980 29474
rect 45461 29416 45466 29472
rect 45522 29416 46980 29472
rect 45461 29414 46980 29416
rect 45461 29411 45527 29414
rect 46974 29412 46980 29414
rect 47044 29474 47050 29476
rect 47209 29474 47275 29477
rect 47044 29472 47275 29474
rect 47044 29416 47214 29472
rect 47270 29416 47275 29472
rect 47044 29414 47275 29416
rect 47044 29412 47050 29414
rect 47209 29411 47275 29414
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 39205 29338 39271 29341
rect 41137 29338 41203 29341
rect 39205 29336 41203 29338
rect 39205 29280 39210 29336
rect 39266 29280 41142 29336
rect 41198 29280 41203 29336
rect 39205 29278 41203 29280
rect 39205 29275 39271 29278
rect 41137 29275 41203 29278
rect 45829 29338 45895 29341
rect 47853 29338 47919 29341
rect 45829 29336 47919 29338
rect 45829 29280 45834 29336
rect 45890 29280 47858 29336
rect 47914 29280 47919 29336
rect 45829 29278 47919 29280
rect 45829 29275 45895 29278
rect 47853 29275 47919 29278
rect 58249 29338 58315 29341
rect 59200 29338 59800 29368
rect 58249 29336 59800 29338
rect 58249 29280 58254 29336
rect 58310 29280 59800 29336
rect 58249 29278 59800 29280
rect 58249 29275 58315 29278
rect 59200 29248 59800 29278
rect 31293 29202 31359 29205
rect 36353 29202 36419 29205
rect 31293 29200 36419 29202
rect 31293 29144 31298 29200
rect 31354 29144 36358 29200
rect 36414 29144 36419 29200
rect 31293 29142 36419 29144
rect 31293 29139 31359 29142
rect 36353 29139 36419 29142
rect 40953 29202 41019 29205
rect 44265 29202 44331 29205
rect 40953 29200 44331 29202
rect 40953 29144 40958 29200
rect 41014 29144 44270 29200
rect 44326 29144 44331 29200
rect 40953 29142 44331 29144
rect 40953 29139 41019 29142
rect 44265 29139 44331 29142
rect 47945 29202 48011 29205
rect 48221 29202 48287 29205
rect 50337 29202 50403 29205
rect 47945 29200 50403 29202
rect 47945 29144 47950 29200
rect 48006 29144 48226 29200
rect 48282 29144 50342 29200
rect 50398 29144 50403 29200
rect 47945 29142 50403 29144
rect 47945 29139 48011 29142
rect 48221 29139 48287 29142
rect 50337 29139 50403 29142
rect 53373 29202 53439 29205
rect 55397 29202 55463 29205
rect 53373 29200 55463 29202
rect 53373 29144 53378 29200
rect 53434 29144 55402 29200
rect 55458 29144 55463 29200
rect 53373 29142 55463 29144
rect 53373 29139 53439 29142
rect 55397 29139 55463 29142
rect 40493 29068 40559 29069
rect 40493 29064 40540 29068
rect 40604 29066 40610 29068
rect 40493 29008 40498 29064
rect 40493 29004 40540 29008
rect 40604 29006 40650 29066
rect 40604 29004 40610 29006
rect 40493 29003 40559 29004
rect 40309 28930 40375 28933
rect 41229 28930 41295 28933
rect 40309 28928 41295 28930
rect 40309 28872 40314 28928
rect 40370 28872 41234 28928
rect 41290 28872 41295 28928
rect 40309 28870 41295 28872
rect 40309 28867 40375 28870
rect 41229 28867 41295 28870
rect 45921 28930 45987 28933
rect 47117 28930 47183 28933
rect 45921 28928 47183 28930
rect 45921 28872 45926 28928
rect 45982 28872 47122 28928
rect 47178 28872 47183 28928
rect 45921 28870 47183 28872
rect 45921 28867 45987 28870
rect 47117 28867 47183 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 40677 28386 40743 28389
rect 41229 28386 41295 28389
rect 41413 28386 41479 28389
rect 40677 28384 41479 28386
rect 40677 28328 40682 28384
rect 40738 28328 41234 28384
rect 41290 28328 41418 28384
rect 41474 28328 41479 28384
rect 40677 28326 41479 28328
rect 40677 28323 40743 28326
rect 41229 28323 41295 28326
rect 41413 28323 41479 28326
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 34329 28252 34395 28253
rect 34278 28188 34284 28252
rect 34348 28250 34395 28252
rect 49601 28250 49667 28253
rect 51993 28250 52059 28253
rect 34348 28248 34440 28250
rect 34390 28192 34440 28248
rect 34348 28190 34440 28192
rect 49601 28248 52059 28250
rect 49601 28192 49606 28248
rect 49662 28192 51998 28248
rect 52054 28192 52059 28248
rect 49601 28190 52059 28192
rect 34348 28188 34395 28190
rect 34329 28187 34395 28188
rect 49601 28187 49667 28190
rect 51993 28187 52059 28190
rect 39481 28114 39547 28117
rect 42517 28114 42583 28117
rect 39481 28112 42583 28114
rect 39481 28056 39486 28112
rect 39542 28056 42522 28112
rect 42578 28056 42583 28112
rect 39481 28054 42583 28056
rect 39481 28051 39547 28054
rect 42517 28051 42583 28054
rect 48957 28114 49023 28117
rect 51073 28114 51139 28117
rect 48957 28112 51139 28114
rect 48957 28056 48962 28112
rect 49018 28056 51078 28112
rect 51134 28056 51139 28112
rect 48957 28054 51139 28056
rect 48957 28051 49023 28054
rect 51073 28051 51139 28054
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 47945 27706 48011 27709
rect 51901 27706 51967 27709
rect 53097 27706 53163 27709
rect 47945 27704 53163 27706
rect 47945 27648 47950 27704
rect 48006 27648 51906 27704
rect 51962 27648 53102 27704
rect 53158 27648 53163 27704
rect 47945 27646 53163 27648
rect 47945 27643 48011 27646
rect 51901 27643 51967 27646
rect 53097 27643 53163 27646
rect 48262 27508 48268 27572
rect 48332 27570 48338 27572
rect 51625 27570 51691 27573
rect 48332 27568 51691 27570
rect 48332 27512 51630 27568
rect 51686 27512 51691 27568
rect 48332 27510 51691 27512
rect 48332 27508 48338 27510
rect 51625 27507 51691 27510
rect 40534 27236 40540 27300
rect 40604 27298 40610 27300
rect 45553 27298 45619 27301
rect 40604 27296 45619 27298
rect 40604 27240 45558 27296
rect 45614 27240 45619 27296
rect 40604 27238 45619 27240
rect 40604 27236 40610 27238
rect 45553 27235 45619 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 35590 27167 35906 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 40125 26618 40191 26621
rect 46657 26618 46723 26621
rect 40125 26616 46723 26618
rect 40125 26560 40130 26616
rect 40186 26560 46662 26616
rect 46718 26560 46723 26616
rect 40125 26558 46723 26560
rect 40125 26555 40191 26558
rect 46657 26555 46723 26558
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 46933 26076 46999 26077
rect 46933 26074 46980 26076
rect 46888 26072 46980 26074
rect 46888 26016 46938 26072
rect 46888 26014 46980 26016
rect 46933 26012 46980 26014
rect 47044 26012 47050 26076
rect 46933 26011 46999 26012
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 39021 24170 39087 24173
rect 41597 24170 41663 24173
rect 39021 24168 41663 24170
rect 39021 24112 39026 24168
rect 39082 24112 41602 24168
rect 41658 24112 41663 24168
rect 39021 24110 41663 24112
rect 39021 24107 39087 24110
rect 41597 24107 41663 24110
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 35590 16287 35906 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
<< via3 >>
rect 4876 57692 4940 57696
rect 4876 57636 4880 57692
rect 4880 57636 4936 57692
rect 4936 57636 4940 57692
rect 4876 57632 4940 57636
rect 4956 57692 5020 57696
rect 4956 57636 4960 57692
rect 4960 57636 5016 57692
rect 5016 57636 5020 57692
rect 4956 57632 5020 57636
rect 5036 57692 5100 57696
rect 5036 57636 5040 57692
rect 5040 57636 5096 57692
rect 5096 57636 5100 57692
rect 5036 57632 5100 57636
rect 5116 57692 5180 57696
rect 5116 57636 5120 57692
rect 5120 57636 5176 57692
rect 5176 57636 5180 57692
rect 5116 57632 5180 57636
rect 35596 57692 35660 57696
rect 35596 57636 35600 57692
rect 35600 57636 35656 57692
rect 35656 57636 35660 57692
rect 35596 57632 35660 57636
rect 35676 57692 35740 57696
rect 35676 57636 35680 57692
rect 35680 57636 35736 57692
rect 35736 57636 35740 57692
rect 35676 57632 35740 57636
rect 35756 57692 35820 57696
rect 35756 57636 35760 57692
rect 35760 57636 35816 57692
rect 35816 57636 35820 57692
rect 35756 57632 35820 57636
rect 35836 57692 35900 57696
rect 35836 57636 35840 57692
rect 35840 57636 35896 57692
rect 35896 57636 35900 57692
rect 35836 57632 35900 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 4876 56604 4940 56608
rect 4876 56548 4880 56604
rect 4880 56548 4936 56604
rect 4936 56548 4940 56604
rect 4876 56544 4940 56548
rect 4956 56604 5020 56608
rect 4956 56548 4960 56604
rect 4960 56548 5016 56604
rect 5016 56548 5020 56604
rect 4956 56544 5020 56548
rect 5036 56604 5100 56608
rect 5036 56548 5040 56604
rect 5040 56548 5096 56604
rect 5096 56548 5100 56604
rect 5036 56544 5100 56548
rect 5116 56604 5180 56608
rect 5116 56548 5120 56604
rect 5120 56548 5176 56604
rect 5176 56548 5180 56604
rect 5116 56544 5180 56548
rect 35596 56604 35660 56608
rect 35596 56548 35600 56604
rect 35600 56548 35656 56604
rect 35656 56548 35660 56604
rect 35596 56544 35660 56548
rect 35676 56604 35740 56608
rect 35676 56548 35680 56604
rect 35680 56548 35736 56604
rect 35736 56548 35740 56604
rect 35676 56544 35740 56548
rect 35756 56604 35820 56608
rect 35756 56548 35760 56604
rect 35760 56548 35816 56604
rect 35816 56548 35820 56604
rect 35756 56544 35820 56548
rect 35836 56604 35900 56608
rect 35836 56548 35840 56604
rect 35840 56548 35896 56604
rect 35896 56548 35900 56604
rect 35836 56544 35900 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 4876 55516 4940 55520
rect 4876 55460 4880 55516
rect 4880 55460 4936 55516
rect 4936 55460 4940 55516
rect 4876 55456 4940 55460
rect 4956 55516 5020 55520
rect 4956 55460 4960 55516
rect 4960 55460 5016 55516
rect 5016 55460 5020 55516
rect 4956 55456 5020 55460
rect 5036 55516 5100 55520
rect 5036 55460 5040 55516
rect 5040 55460 5096 55516
rect 5096 55460 5100 55516
rect 5036 55456 5100 55460
rect 5116 55516 5180 55520
rect 5116 55460 5120 55516
rect 5120 55460 5176 55516
rect 5176 55460 5180 55516
rect 5116 55456 5180 55460
rect 35596 55516 35660 55520
rect 35596 55460 35600 55516
rect 35600 55460 35656 55516
rect 35656 55460 35660 55516
rect 35596 55456 35660 55460
rect 35676 55516 35740 55520
rect 35676 55460 35680 55516
rect 35680 55460 35736 55516
rect 35736 55460 35740 55516
rect 35676 55456 35740 55460
rect 35756 55516 35820 55520
rect 35756 55460 35760 55516
rect 35760 55460 35816 55516
rect 35816 55460 35820 55516
rect 35756 55456 35820 55460
rect 35836 55516 35900 55520
rect 35836 55460 35840 55516
rect 35840 55460 35896 55516
rect 35896 55460 35900 55516
rect 35836 55456 35900 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 4876 54428 4940 54432
rect 4876 54372 4880 54428
rect 4880 54372 4936 54428
rect 4936 54372 4940 54428
rect 4876 54368 4940 54372
rect 4956 54428 5020 54432
rect 4956 54372 4960 54428
rect 4960 54372 5016 54428
rect 5016 54372 5020 54428
rect 4956 54368 5020 54372
rect 5036 54428 5100 54432
rect 5036 54372 5040 54428
rect 5040 54372 5096 54428
rect 5096 54372 5100 54428
rect 5036 54368 5100 54372
rect 5116 54428 5180 54432
rect 5116 54372 5120 54428
rect 5120 54372 5176 54428
rect 5176 54372 5180 54428
rect 5116 54368 5180 54372
rect 35596 54428 35660 54432
rect 35596 54372 35600 54428
rect 35600 54372 35656 54428
rect 35656 54372 35660 54428
rect 35596 54368 35660 54372
rect 35676 54428 35740 54432
rect 35676 54372 35680 54428
rect 35680 54372 35736 54428
rect 35736 54372 35740 54428
rect 35676 54368 35740 54372
rect 35756 54428 35820 54432
rect 35756 54372 35760 54428
rect 35760 54372 35816 54428
rect 35816 54372 35820 54428
rect 35756 54368 35820 54372
rect 35836 54428 35900 54432
rect 35836 54372 35840 54428
rect 35840 54372 35896 54428
rect 35896 54372 35900 54428
rect 35836 54368 35900 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 4876 53340 4940 53344
rect 4876 53284 4880 53340
rect 4880 53284 4936 53340
rect 4936 53284 4940 53340
rect 4876 53280 4940 53284
rect 4956 53340 5020 53344
rect 4956 53284 4960 53340
rect 4960 53284 5016 53340
rect 5016 53284 5020 53340
rect 4956 53280 5020 53284
rect 5036 53340 5100 53344
rect 5036 53284 5040 53340
rect 5040 53284 5096 53340
rect 5096 53284 5100 53340
rect 5036 53280 5100 53284
rect 5116 53340 5180 53344
rect 5116 53284 5120 53340
rect 5120 53284 5176 53340
rect 5176 53284 5180 53340
rect 5116 53280 5180 53284
rect 35596 53340 35660 53344
rect 35596 53284 35600 53340
rect 35600 53284 35656 53340
rect 35656 53284 35660 53340
rect 35596 53280 35660 53284
rect 35676 53340 35740 53344
rect 35676 53284 35680 53340
rect 35680 53284 35736 53340
rect 35736 53284 35740 53340
rect 35676 53280 35740 53284
rect 35756 53340 35820 53344
rect 35756 53284 35760 53340
rect 35760 53284 35816 53340
rect 35816 53284 35820 53340
rect 35756 53280 35820 53284
rect 35836 53340 35900 53344
rect 35836 53284 35840 53340
rect 35840 53284 35896 53340
rect 35896 53284 35900 53340
rect 35836 53280 35900 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 4876 52252 4940 52256
rect 4876 52196 4880 52252
rect 4880 52196 4936 52252
rect 4936 52196 4940 52252
rect 4876 52192 4940 52196
rect 4956 52252 5020 52256
rect 4956 52196 4960 52252
rect 4960 52196 5016 52252
rect 5016 52196 5020 52252
rect 4956 52192 5020 52196
rect 5036 52252 5100 52256
rect 5036 52196 5040 52252
rect 5040 52196 5096 52252
rect 5096 52196 5100 52252
rect 5036 52192 5100 52196
rect 5116 52252 5180 52256
rect 5116 52196 5120 52252
rect 5120 52196 5176 52252
rect 5176 52196 5180 52252
rect 5116 52192 5180 52196
rect 35596 52252 35660 52256
rect 35596 52196 35600 52252
rect 35600 52196 35656 52252
rect 35656 52196 35660 52252
rect 35596 52192 35660 52196
rect 35676 52252 35740 52256
rect 35676 52196 35680 52252
rect 35680 52196 35736 52252
rect 35736 52196 35740 52252
rect 35676 52192 35740 52196
rect 35756 52252 35820 52256
rect 35756 52196 35760 52252
rect 35760 52196 35816 52252
rect 35816 52196 35820 52252
rect 35756 52192 35820 52196
rect 35836 52252 35900 52256
rect 35836 52196 35840 52252
rect 35840 52196 35896 52252
rect 35896 52196 35900 52252
rect 35836 52192 35900 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 4876 51164 4940 51168
rect 4876 51108 4880 51164
rect 4880 51108 4936 51164
rect 4936 51108 4940 51164
rect 4876 51104 4940 51108
rect 4956 51164 5020 51168
rect 4956 51108 4960 51164
rect 4960 51108 5016 51164
rect 5016 51108 5020 51164
rect 4956 51104 5020 51108
rect 5036 51164 5100 51168
rect 5036 51108 5040 51164
rect 5040 51108 5096 51164
rect 5096 51108 5100 51164
rect 5036 51104 5100 51108
rect 5116 51164 5180 51168
rect 5116 51108 5120 51164
rect 5120 51108 5176 51164
rect 5176 51108 5180 51164
rect 5116 51104 5180 51108
rect 35596 51164 35660 51168
rect 35596 51108 35600 51164
rect 35600 51108 35656 51164
rect 35656 51108 35660 51164
rect 35596 51104 35660 51108
rect 35676 51164 35740 51168
rect 35676 51108 35680 51164
rect 35680 51108 35736 51164
rect 35736 51108 35740 51164
rect 35676 51104 35740 51108
rect 35756 51164 35820 51168
rect 35756 51108 35760 51164
rect 35760 51108 35816 51164
rect 35816 51108 35820 51164
rect 35756 51104 35820 51108
rect 35836 51164 35900 51168
rect 35836 51108 35840 51164
rect 35840 51108 35896 51164
rect 35896 51108 35900 51164
rect 35836 51104 35900 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 4876 50076 4940 50080
rect 4876 50020 4880 50076
rect 4880 50020 4936 50076
rect 4936 50020 4940 50076
rect 4876 50016 4940 50020
rect 4956 50076 5020 50080
rect 4956 50020 4960 50076
rect 4960 50020 5016 50076
rect 5016 50020 5020 50076
rect 4956 50016 5020 50020
rect 5036 50076 5100 50080
rect 5036 50020 5040 50076
rect 5040 50020 5096 50076
rect 5096 50020 5100 50076
rect 5036 50016 5100 50020
rect 5116 50076 5180 50080
rect 5116 50020 5120 50076
rect 5120 50020 5176 50076
rect 5176 50020 5180 50076
rect 5116 50016 5180 50020
rect 35596 50076 35660 50080
rect 35596 50020 35600 50076
rect 35600 50020 35656 50076
rect 35656 50020 35660 50076
rect 35596 50016 35660 50020
rect 35676 50076 35740 50080
rect 35676 50020 35680 50076
rect 35680 50020 35736 50076
rect 35736 50020 35740 50076
rect 35676 50016 35740 50020
rect 35756 50076 35820 50080
rect 35756 50020 35760 50076
rect 35760 50020 35816 50076
rect 35816 50020 35820 50076
rect 35756 50016 35820 50020
rect 35836 50076 35900 50080
rect 35836 50020 35840 50076
rect 35840 50020 35896 50076
rect 35896 50020 35900 50076
rect 35836 50016 35900 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 4876 48988 4940 48992
rect 4876 48932 4880 48988
rect 4880 48932 4936 48988
rect 4936 48932 4940 48988
rect 4876 48928 4940 48932
rect 4956 48988 5020 48992
rect 4956 48932 4960 48988
rect 4960 48932 5016 48988
rect 5016 48932 5020 48988
rect 4956 48928 5020 48932
rect 5036 48988 5100 48992
rect 5036 48932 5040 48988
rect 5040 48932 5096 48988
rect 5096 48932 5100 48988
rect 5036 48928 5100 48932
rect 5116 48988 5180 48992
rect 5116 48932 5120 48988
rect 5120 48932 5176 48988
rect 5176 48932 5180 48988
rect 5116 48928 5180 48932
rect 35596 48988 35660 48992
rect 35596 48932 35600 48988
rect 35600 48932 35656 48988
rect 35656 48932 35660 48988
rect 35596 48928 35660 48932
rect 35676 48988 35740 48992
rect 35676 48932 35680 48988
rect 35680 48932 35736 48988
rect 35736 48932 35740 48988
rect 35676 48928 35740 48932
rect 35756 48988 35820 48992
rect 35756 48932 35760 48988
rect 35760 48932 35816 48988
rect 35816 48932 35820 48988
rect 35756 48928 35820 48932
rect 35836 48988 35900 48992
rect 35836 48932 35840 48988
rect 35840 48932 35896 48988
rect 35896 48932 35900 48988
rect 35836 48928 35900 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 4876 47900 4940 47904
rect 4876 47844 4880 47900
rect 4880 47844 4936 47900
rect 4936 47844 4940 47900
rect 4876 47840 4940 47844
rect 4956 47900 5020 47904
rect 4956 47844 4960 47900
rect 4960 47844 5016 47900
rect 5016 47844 5020 47900
rect 4956 47840 5020 47844
rect 5036 47900 5100 47904
rect 5036 47844 5040 47900
rect 5040 47844 5096 47900
rect 5096 47844 5100 47900
rect 5036 47840 5100 47844
rect 5116 47900 5180 47904
rect 5116 47844 5120 47900
rect 5120 47844 5176 47900
rect 5176 47844 5180 47900
rect 5116 47840 5180 47844
rect 35596 47900 35660 47904
rect 35596 47844 35600 47900
rect 35600 47844 35656 47900
rect 35656 47844 35660 47900
rect 35596 47840 35660 47844
rect 35676 47900 35740 47904
rect 35676 47844 35680 47900
rect 35680 47844 35736 47900
rect 35736 47844 35740 47900
rect 35676 47840 35740 47844
rect 35756 47900 35820 47904
rect 35756 47844 35760 47900
rect 35760 47844 35816 47900
rect 35816 47844 35820 47900
rect 35756 47840 35820 47844
rect 35836 47900 35900 47904
rect 35836 47844 35840 47900
rect 35840 47844 35896 47900
rect 35896 47844 35900 47900
rect 35836 47840 35900 47844
rect 42012 47364 42076 47428
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 4876 46812 4940 46816
rect 4876 46756 4880 46812
rect 4880 46756 4936 46812
rect 4936 46756 4940 46812
rect 4876 46752 4940 46756
rect 4956 46812 5020 46816
rect 4956 46756 4960 46812
rect 4960 46756 5016 46812
rect 5016 46756 5020 46812
rect 4956 46752 5020 46756
rect 5036 46812 5100 46816
rect 5036 46756 5040 46812
rect 5040 46756 5096 46812
rect 5096 46756 5100 46812
rect 5036 46752 5100 46756
rect 5116 46812 5180 46816
rect 5116 46756 5120 46812
rect 5120 46756 5176 46812
rect 5176 46756 5180 46812
rect 5116 46752 5180 46756
rect 35596 46812 35660 46816
rect 35596 46756 35600 46812
rect 35600 46756 35656 46812
rect 35656 46756 35660 46812
rect 35596 46752 35660 46756
rect 35676 46812 35740 46816
rect 35676 46756 35680 46812
rect 35680 46756 35736 46812
rect 35736 46756 35740 46812
rect 35676 46752 35740 46756
rect 35756 46812 35820 46816
rect 35756 46756 35760 46812
rect 35760 46756 35816 46812
rect 35816 46756 35820 46812
rect 35756 46752 35820 46756
rect 35836 46812 35900 46816
rect 35836 46756 35840 46812
rect 35840 46756 35896 46812
rect 35896 46756 35900 46812
rect 35836 46752 35900 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 42012 45868 42076 45932
rect 32444 45732 32508 45796
rect 4876 45724 4940 45728
rect 4876 45668 4880 45724
rect 4880 45668 4936 45724
rect 4936 45668 4940 45724
rect 4876 45664 4940 45668
rect 4956 45724 5020 45728
rect 4956 45668 4960 45724
rect 4960 45668 5016 45724
rect 5016 45668 5020 45724
rect 4956 45664 5020 45668
rect 5036 45724 5100 45728
rect 5036 45668 5040 45724
rect 5040 45668 5096 45724
rect 5096 45668 5100 45724
rect 5036 45664 5100 45668
rect 5116 45724 5180 45728
rect 5116 45668 5120 45724
rect 5120 45668 5176 45724
rect 5176 45668 5180 45724
rect 5116 45664 5180 45668
rect 35596 45724 35660 45728
rect 35596 45668 35600 45724
rect 35600 45668 35656 45724
rect 35656 45668 35660 45724
rect 35596 45664 35660 45668
rect 35676 45724 35740 45728
rect 35676 45668 35680 45724
rect 35680 45668 35736 45724
rect 35736 45668 35740 45724
rect 35676 45664 35740 45668
rect 35756 45724 35820 45728
rect 35756 45668 35760 45724
rect 35760 45668 35816 45724
rect 35816 45668 35820 45724
rect 35756 45664 35820 45668
rect 35836 45724 35900 45728
rect 35836 45668 35840 45724
rect 35840 45668 35896 45724
rect 35896 45668 35900 45724
rect 35836 45664 35900 45668
rect 48636 45596 48700 45660
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 37596 44780 37660 44844
rect 4876 44636 4940 44640
rect 4876 44580 4880 44636
rect 4880 44580 4936 44636
rect 4936 44580 4940 44636
rect 4876 44576 4940 44580
rect 4956 44636 5020 44640
rect 4956 44580 4960 44636
rect 4960 44580 5016 44636
rect 5016 44580 5020 44636
rect 4956 44576 5020 44580
rect 5036 44636 5100 44640
rect 5036 44580 5040 44636
rect 5040 44580 5096 44636
rect 5096 44580 5100 44636
rect 5036 44576 5100 44580
rect 5116 44636 5180 44640
rect 5116 44580 5120 44636
rect 5120 44580 5176 44636
rect 5176 44580 5180 44636
rect 5116 44576 5180 44580
rect 35596 44636 35660 44640
rect 35596 44580 35600 44636
rect 35600 44580 35656 44636
rect 35656 44580 35660 44636
rect 35596 44576 35660 44580
rect 35676 44636 35740 44640
rect 35676 44580 35680 44636
rect 35680 44580 35736 44636
rect 35736 44580 35740 44636
rect 35676 44576 35740 44580
rect 35756 44636 35820 44640
rect 35756 44580 35760 44636
rect 35760 44580 35816 44636
rect 35816 44580 35820 44636
rect 35756 44576 35820 44580
rect 35836 44636 35900 44640
rect 35836 44580 35840 44636
rect 35840 44580 35896 44636
rect 35896 44580 35900 44636
rect 35836 44576 35900 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 35596 43548 35660 43552
rect 35596 43492 35600 43548
rect 35600 43492 35656 43548
rect 35656 43492 35660 43548
rect 35596 43488 35660 43492
rect 35676 43548 35740 43552
rect 35676 43492 35680 43548
rect 35680 43492 35736 43548
rect 35736 43492 35740 43548
rect 35676 43488 35740 43492
rect 35756 43548 35820 43552
rect 35756 43492 35760 43548
rect 35760 43492 35816 43548
rect 35816 43492 35820 43548
rect 35756 43488 35820 43492
rect 35836 43548 35900 43552
rect 35836 43492 35840 43548
rect 35840 43492 35896 43548
rect 35896 43492 35900 43548
rect 35836 43488 35900 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 41092 42876 41156 42940
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 35596 42460 35660 42464
rect 35596 42404 35600 42460
rect 35600 42404 35656 42460
rect 35656 42404 35660 42460
rect 35596 42400 35660 42404
rect 35676 42460 35740 42464
rect 35676 42404 35680 42460
rect 35680 42404 35736 42460
rect 35736 42404 35740 42460
rect 35676 42400 35740 42404
rect 35756 42460 35820 42464
rect 35756 42404 35760 42460
rect 35760 42404 35816 42460
rect 35816 42404 35820 42460
rect 35756 42400 35820 42404
rect 35836 42460 35900 42464
rect 35836 42404 35840 42460
rect 35840 42404 35896 42460
rect 35896 42404 35900 42460
rect 35836 42400 35900 42404
rect 34284 41924 34348 41988
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 35596 41372 35660 41376
rect 35596 41316 35600 41372
rect 35600 41316 35656 41372
rect 35656 41316 35660 41372
rect 35596 41312 35660 41316
rect 35676 41372 35740 41376
rect 35676 41316 35680 41372
rect 35680 41316 35736 41372
rect 35736 41316 35740 41372
rect 35676 41312 35740 41316
rect 35756 41372 35820 41376
rect 35756 41316 35760 41372
rect 35760 41316 35816 41372
rect 35816 41316 35820 41372
rect 35756 41312 35820 41316
rect 35836 41372 35900 41376
rect 35836 41316 35840 41372
rect 35840 41316 35896 41372
rect 35896 41316 35900 41372
rect 35836 41312 35900 41316
rect 38516 41304 38580 41308
rect 38516 41248 38566 41304
rect 38566 41248 38580 41304
rect 38516 41244 38580 41248
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 38516 40700 38580 40764
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 35596 40284 35660 40288
rect 35596 40228 35600 40284
rect 35600 40228 35656 40284
rect 35656 40228 35660 40284
rect 35596 40224 35660 40228
rect 35676 40284 35740 40288
rect 35676 40228 35680 40284
rect 35680 40228 35736 40284
rect 35736 40228 35740 40284
rect 35676 40224 35740 40228
rect 35756 40284 35820 40288
rect 35756 40228 35760 40284
rect 35760 40228 35816 40284
rect 35816 40228 35820 40284
rect 35756 40224 35820 40228
rect 35836 40284 35900 40288
rect 35836 40228 35840 40284
rect 35840 40228 35896 40284
rect 35896 40228 35900 40284
rect 35836 40224 35900 40228
rect 48268 39944 48332 39948
rect 48268 39888 48318 39944
rect 48318 39888 48332 39944
rect 48268 39884 48332 39888
rect 48636 39884 48700 39948
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 35596 39196 35660 39200
rect 35596 39140 35600 39196
rect 35600 39140 35656 39196
rect 35656 39140 35660 39196
rect 35596 39136 35660 39140
rect 35676 39196 35740 39200
rect 35676 39140 35680 39196
rect 35680 39140 35736 39196
rect 35736 39140 35740 39196
rect 35676 39136 35740 39140
rect 35756 39196 35820 39200
rect 35756 39140 35760 39196
rect 35760 39140 35816 39196
rect 35816 39140 35820 39196
rect 35756 39136 35820 39140
rect 35836 39196 35900 39200
rect 35836 39140 35840 39196
rect 35840 39140 35896 39196
rect 35896 39140 35900 39196
rect 35836 39136 35900 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 35596 38108 35660 38112
rect 35596 38052 35600 38108
rect 35600 38052 35656 38108
rect 35656 38052 35660 38108
rect 35596 38048 35660 38052
rect 35676 38108 35740 38112
rect 35676 38052 35680 38108
rect 35680 38052 35736 38108
rect 35736 38052 35740 38108
rect 35676 38048 35740 38052
rect 35756 38108 35820 38112
rect 35756 38052 35760 38108
rect 35760 38052 35816 38108
rect 35816 38052 35820 38108
rect 35756 38048 35820 38052
rect 35836 38108 35900 38112
rect 35836 38052 35840 38108
rect 35840 38052 35896 38108
rect 35896 38052 35900 38108
rect 35836 38048 35900 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 42012 33084 42076 33148
rect 48268 33084 48332 33148
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 37596 32600 37660 32604
rect 37596 32544 37610 32600
rect 37610 32544 37660 32600
rect 37596 32540 37660 32544
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 41092 31860 41156 31924
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 48268 30364 48332 30428
rect 32444 30288 32508 30292
rect 32444 30232 32458 30288
rect 32458 30232 32508 30288
rect 32444 30228 32508 30232
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 46980 29412 47044 29476
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 40540 29064 40604 29068
rect 40540 29008 40554 29064
rect 40554 29008 40604 29064
rect 40540 29004 40604 29008
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 34284 28248 34348 28252
rect 34284 28192 34334 28248
rect 34334 28192 34348 28248
rect 34284 28188 34348 28192
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 48268 27508 48332 27572
rect 40540 27236 40604 27300
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 46980 26072 47044 26076
rect 46980 26016 46994 26072
rect 46994 26016 47044 26072
rect 46980 26012 47044 26016
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 57696 5188 57712
rect 4868 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5188 57696
rect 4868 56608 5188 57632
rect 4868 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5188 56608
rect 4868 55520 5188 56544
rect 4868 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5188 55520
rect 4868 54432 5188 55456
rect 4868 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5188 54432
rect 4868 53344 5188 54368
rect 4868 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5188 53344
rect 4868 52256 5188 53280
rect 4868 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5188 52256
rect 4868 51168 5188 52192
rect 4868 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5188 51168
rect 4868 50080 5188 51104
rect 4868 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5188 50080
rect 4868 48992 5188 50016
rect 4868 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5188 48992
rect 4868 47904 5188 48928
rect 4868 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5188 47904
rect 4868 46816 5188 47840
rect 4868 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5188 46816
rect 4868 45728 5188 46752
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 32443 45796 32509 45797
rect 32443 45732 32444 45796
rect 32508 45732 32509 45796
rect 32443 45731 32509 45732
rect 4868 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5188 45728
rect 4868 44640 5188 45664
rect 4868 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5188 44640
rect 4868 43552 5188 44576
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 32446 30293 32506 45731
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34283 41988 34349 41989
rect 34283 41924 34284 41988
rect 34348 41924 34349 41988
rect 34283 41923 34349 41924
rect 32443 30292 32509 30293
rect 32443 30228 32444 30292
rect 32508 30228 32509 30292
rect 32443 30227 32509 30228
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 34286 28253 34346 41923
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36260 35248 36416
rect 34928 36024 34970 36260
rect 35206 36024 35248 36260
rect 34928 35392 35248 36024
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34283 28252 34349 28253
rect 34283 28188 34284 28252
rect 34348 28188 34349 28252
rect 34283 28187 34349 28188
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 57696 35908 57712
rect 35588 57632 35596 57696
rect 35660 57632 35676 57696
rect 35740 57632 35756 57696
rect 35820 57632 35836 57696
rect 35900 57632 35908 57696
rect 35588 56608 35908 57632
rect 35588 56544 35596 56608
rect 35660 56544 35676 56608
rect 35740 56544 35756 56608
rect 35820 56544 35836 56608
rect 35900 56544 35908 56608
rect 35588 55520 35908 56544
rect 35588 55456 35596 55520
rect 35660 55456 35676 55520
rect 35740 55456 35756 55520
rect 35820 55456 35836 55520
rect 35900 55456 35908 55520
rect 35588 54432 35908 55456
rect 35588 54368 35596 54432
rect 35660 54368 35676 54432
rect 35740 54368 35756 54432
rect 35820 54368 35836 54432
rect 35900 54368 35908 54432
rect 35588 53344 35908 54368
rect 35588 53280 35596 53344
rect 35660 53280 35676 53344
rect 35740 53280 35756 53344
rect 35820 53280 35836 53344
rect 35900 53280 35908 53344
rect 35588 52256 35908 53280
rect 35588 52192 35596 52256
rect 35660 52192 35676 52256
rect 35740 52192 35756 52256
rect 35820 52192 35836 52256
rect 35900 52192 35908 52256
rect 35588 51168 35908 52192
rect 35588 51104 35596 51168
rect 35660 51104 35676 51168
rect 35740 51104 35756 51168
rect 35820 51104 35836 51168
rect 35900 51104 35908 51168
rect 35588 50080 35908 51104
rect 35588 50016 35596 50080
rect 35660 50016 35676 50080
rect 35740 50016 35756 50080
rect 35820 50016 35836 50080
rect 35900 50016 35908 50080
rect 35588 48992 35908 50016
rect 35588 48928 35596 48992
rect 35660 48928 35676 48992
rect 35740 48928 35756 48992
rect 35820 48928 35836 48992
rect 35900 48928 35908 48992
rect 35588 47904 35908 48928
rect 35588 47840 35596 47904
rect 35660 47840 35676 47904
rect 35740 47840 35756 47904
rect 35820 47840 35836 47904
rect 35900 47840 35908 47904
rect 35588 46816 35908 47840
rect 42011 47428 42077 47429
rect 42011 47364 42012 47428
rect 42076 47364 42077 47428
rect 42011 47363 42077 47364
rect 35588 46752 35596 46816
rect 35660 46752 35676 46816
rect 35740 46752 35756 46816
rect 35820 46752 35836 46816
rect 35900 46752 35908 46816
rect 35588 45728 35908 46752
rect 42014 45933 42074 47363
rect 42011 45932 42077 45933
rect 42011 45868 42012 45932
rect 42076 45868 42077 45932
rect 42011 45867 42077 45868
rect 35588 45664 35596 45728
rect 35660 45664 35676 45728
rect 35740 45664 35756 45728
rect 35820 45664 35836 45728
rect 35900 45664 35908 45728
rect 35588 44640 35908 45664
rect 37595 44844 37661 44845
rect 37595 44780 37596 44844
rect 37660 44780 37661 44844
rect 37595 44779 37661 44780
rect 35588 44576 35596 44640
rect 35660 44576 35676 44640
rect 35740 44576 35756 44640
rect 35820 44576 35836 44640
rect 35900 44576 35908 44640
rect 35588 43552 35908 44576
rect 35588 43488 35596 43552
rect 35660 43488 35676 43552
rect 35740 43488 35756 43552
rect 35820 43488 35836 43552
rect 35900 43488 35908 43552
rect 35588 42464 35908 43488
rect 35588 42400 35596 42464
rect 35660 42400 35676 42464
rect 35740 42400 35756 42464
rect 35820 42400 35836 42464
rect 35900 42400 35908 42464
rect 35588 41376 35908 42400
rect 35588 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35908 41376
rect 35588 40288 35908 41312
rect 35588 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35908 40288
rect 35588 39200 35908 40224
rect 35588 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35908 39200
rect 35588 38112 35908 39136
rect 35588 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35908 38112
rect 35588 37024 35908 38048
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 36920 35908 36960
rect 35588 36684 35630 36920
rect 35866 36684 35908 36920
rect 35588 35936 35908 36684
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 37598 32605 37658 44779
rect 41091 42940 41157 42941
rect 41091 42876 41092 42940
rect 41156 42876 41157 42940
rect 41091 42875 41157 42876
rect 38515 41308 38581 41309
rect 38515 41244 38516 41308
rect 38580 41244 38581 41308
rect 38515 41243 38581 41244
rect 38518 40765 38578 41243
rect 38515 40764 38581 40765
rect 38515 40700 38516 40764
rect 38580 40700 38581 40764
rect 38515 40699 38581 40700
rect 37595 32604 37661 32605
rect 37595 32540 37596 32604
rect 37660 32540 37661 32604
rect 37595 32539 37661 32540
rect 41094 31925 41154 42875
rect 42014 33149 42074 45867
rect 48635 45660 48701 45661
rect 48635 45596 48636 45660
rect 48700 45596 48701 45660
rect 48635 45595 48701 45596
rect 48638 39949 48698 45595
rect 48267 39948 48333 39949
rect 48267 39884 48268 39948
rect 48332 39884 48333 39948
rect 48267 39883 48333 39884
rect 48635 39948 48701 39949
rect 48635 39884 48636 39948
rect 48700 39884 48701 39948
rect 48635 39883 48701 39884
rect 48270 33149 48330 39883
rect 42011 33148 42077 33149
rect 42011 33084 42012 33148
rect 42076 33084 42077 33148
rect 42011 33083 42077 33084
rect 48267 33148 48333 33149
rect 48267 33084 48268 33148
rect 48332 33084 48333 33148
rect 48267 33083 48333 33084
rect 41091 31924 41157 31925
rect 41091 31860 41092 31924
rect 41156 31860 41157 31924
rect 41091 31859 41157 31860
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 48267 30428 48333 30429
rect 48267 30364 48268 30428
rect 48332 30364 48333 30428
rect 48267 30363 48333 30364
rect 46979 29476 47045 29477
rect 46979 29412 46980 29476
rect 47044 29412 47045 29476
rect 46979 29411 47045 29412
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 40539 29068 40605 29069
rect 40539 29004 40540 29068
rect 40604 29004 40605 29068
rect 40539 29003 40605 29004
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 40542 27301 40602 29003
rect 40539 27300 40605 27301
rect 40539 27236 40540 27300
rect 40604 27236 40605 27300
rect 40539 27235 40605 27236
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 46982 26077 47042 29411
rect 48270 27573 48330 30363
rect 48267 27572 48333 27573
rect 48267 27508 48268 27572
rect 48332 27508 48333 27572
rect 48267 27507 48333 27508
rect 46979 26076 47045 26077
rect 46979 26012 46980 26076
rect 47044 26012 47045 26076
rect 46979 26011 47045 26012
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
<< via4 >>
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 36684 5146 36920
rect 34970 36024 35206 36260
rect 4910 6048 5146 6284
rect 34970 5388 35206 5624
rect 35630 36684 35866 36920
rect 35630 6048 35866 6284
<< metal5 >>
rect 1056 36920 58928 36962
rect 1056 36684 4910 36920
rect 5146 36684 35630 36920
rect 35866 36684 58928 36920
rect 1056 36642 58928 36684
rect 1056 36260 58928 36302
rect 1056 36024 4250 36260
rect 4486 36024 34970 36260
rect 35206 36024 58928 36260
rect 1056 35982 58928 36024
rect 1056 6284 58928 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 58928 6284
rect 1056 6006 58928 6048
rect 1056 5624 58928 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 58928 5624
rect 1056 5346 58928 5388
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A0 OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 47288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A
timestamp 1667941163
transform 1 0 57316 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A
timestamp 1667941163
transform -1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A1
timestamp 1667941163
transform 1 0 49588 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A
timestamp 1667941163
transform 1 0 33672 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A
timestamp 1667941163
transform -1 0 42780 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A1
timestamp 1667941163
transform 1 0 41308 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A
timestamp 1667941163
transform -1 0 39468 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A0
timestamp 1667941163
transform 1 0 36800 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A1
timestamp 1667941163
transform 1 0 36708 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A1
timestamp 1667941163
transform 1 0 35512 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A1
timestamp 1667941163
transform 1 0 34868 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A
timestamp 1667941163
transform -1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B2
timestamp 1667941163
transform -1 0 44712 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A
timestamp 1667941163
transform 1 0 43240 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__B2
timestamp 1667941163
transform 1 0 47104 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A0
timestamp 1667941163
transform -1 0 43608 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A1
timestamp 1667941163
transform -1 0 44160 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A
timestamp 1667941163
transform 1 0 42596 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A1
timestamp 1667941163
transform 1 0 42136 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__B2
timestamp 1667941163
transform 1 0 45448 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__B2
timestamp 1667941163
transform 1 0 43608 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A
timestamp 1667941163
transform -1 0 33028 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A
timestamp 1667941163
transform 1 0 35604 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A0
timestamp 1667941163
transform -1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A1
timestamp 1667941163
transform -1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A0
timestamp 1667941163
transform 1 0 37628 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A1
timestamp 1667941163
transform 1 0 38180 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1667941163
transform -1 0 33856 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__B2
timestamp 1667941163
transform 1 0 38088 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A
timestamp 1667941163
transform -1 0 42228 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__B2
timestamp 1667941163
transform 1 0 41032 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1667941163
transform -1 0 43608 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A0
timestamp 1667941163
transform -1 0 37628 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A1
timestamp 1667941163
transform 1 0 38180 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A
timestamp 1667941163
transform 1 0 46184 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A1
timestamp 1667941163
transform 1 0 41584 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A
timestamp 1667941163
transform -1 0 47840 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__B2
timestamp 1667941163
transform -1 0 36984 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__B2
timestamp 1667941163
transform 1 0 38732 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A0
timestamp 1667941163
transform 1 0 44896 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A1
timestamp 1667941163
transform -1 0 44712 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A1
timestamp 1667941163
transform 1 0 2392 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__S
timestamp 1667941163
transform -1 0 2944 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1667941163
transform 1 0 51612 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A
timestamp 1667941163
transform 1 0 30728 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A
timestamp 1667941163
transform -1 0 28796 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1667941163
transform 1 0 30360 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A
timestamp 1667941163
transform -1 0 45356 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1667941163
transform 1 0 34224 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A
timestamp 1667941163
transform 1 0 29072 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A
timestamp 1667941163
transform 1 0 31648 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A
timestamp 1667941163
transform 1 0 31464 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__B2
timestamp 1667941163
transform 1 0 40020 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A1
timestamp 1667941163
transform -1 0 39928 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__B2
timestamp 1667941163
transform 1 0 41860 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B1
timestamp 1667941163
transform 1 0 35880 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A1
timestamp 1667941163
transform -1 0 37628 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__B1
timestamp 1667941163
transform -1 0 35512 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__B1
timestamp 1667941163
transform 1 0 39008 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__B1
timestamp 1667941163
transform 1 0 37996 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A1
timestamp 1667941163
transform 1 0 39376 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__B2
timestamp 1667941163
transform 1 0 39008 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__B1
timestamp 1667941163
transform 1 0 37444 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__B1
timestamp 1667941163
transform -1 0 40204 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__B2
timestamp 1667941163
transform 1 0 40572 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A1
timestamp 1667941163
transform 1 0 42596 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A1
timestamp 1667941163
transform 1 0 41400 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A1
timestamp 1667941163
transform -1 0 39468 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__B1
timestamp 1667941163
transform -1 0 36156 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A1
timestamp 1667941163
transform -1 0 36800 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__B1
timestamp 1667941163
transform -1 0 34408 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__S
timestamp 1667941163
transform 1 0 47840 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__B2
timestamp 1667941163
transform -1 0 45356 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__B2
timestamp 1667941163
transform -1 0 41676 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__B1
timestamp 1667941163
transform 1 0 30452 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__A1
timestamp 1667941163
transform -1 0 35052 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__B1
timestamp 1667941163
transform 1 0 34040 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A1
timestamp 1667941163
transform 1 0 33396 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A1
timestamp 1667941163
transform -1 0 31096 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__B1
timestamp 1667941163
transform 1 0 31648 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__B1
timestamp 1667941163
transform -1 0 31280 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__B2
timestamp 1667941163
transform -1 0 34960 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A1
timestamp 1667941163
transform 1 0 33028 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__A1
timestamp 1667941163
transform -1 0 37076 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__B2
timestamp 1667941163
transform -1 0 41952 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__B1
timestamp 1667941163
transform 1 0 45172 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A1
timestamp 1667941163
transform 1 0 45172 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A1
timestamp 1667941163
transform 1 0 44436 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A1
timestamp 1667941163
transform -1 0 44160 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__B2
timestamp 1667941163
transform -1 0 44712 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A
timestamp 1667941163
transform 1 0 52256 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A1
timestamp 1667941163
transform 1 0 49588 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A1
timestamp 1667941163
transform 1 0 33212 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__B2
timestamp 1667941163
transform 1 0 34132 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__B1
timestamp 1667941163
transform -1 0 28796 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A1
timestamp 1667941163
transform 1 0 33120 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__A1
timestamp 1667941163
transform -1 0 44160 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A1
timestamp 1667941163
transform 1 0 41124 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A1
timestamp 1667941163
transform 1 0 34040 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__A1
timestamp 1667941163
transform 1 0 34868 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__B2
timestamp 1667941163
transform 1 0 47104 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A1
timestamp 1667941163
transform 1 0 46276 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__A1
timestamp 1667941163
transform 1 0 49220 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__B2
timestamp 1667941163
transform 1 0 35512 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__B2
timestamp 1667941163
transform -1 0 49404 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__B1
timestamp 1667941163
transform 1 0 47380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A1
timestamp 1667941163
transform -1 0 55384 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__B2
timestamp 1667941163
transform 1 0 46276 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__B2
timestamp 1667941163
transform -1 0 44712 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A1
timestamp 1667941163
transform 1 0 50140 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__B2
timestamp 1667941163
transform 1 0 47564 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__C1
timestamp 1667941163
transform 1 0 52164 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__B1
timestamp 1667941163
transform 1 0 36708 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__A1
timestamp 1667941163
transform 1 0 40020 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__B2
timestamp 1667941163
transform 1 0 40572 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A1
timestamp 1667941163
transform -1 0 36432 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__B1
timestamp 1667941163
transform -1 0 39468 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__B1
timestamp 1667941163
transform 1 0 38180 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__B2
timestamp 1667941163
transform 1 0 39744 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__B
timestamp 1667941163
transform 1 0 50876 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__B1
timestamp 1667941163
transform -1 0 37260 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__A1
timestamp 1667941163
transform 1 0 38548 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__A1
timestamp 1667941163
transform 1 0 38548 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__B1
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1
timestamp 1667941163
transform 1 0 43516 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__B1
timestamp 1667941163
transform 1 0 35604 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__B2
timestamp 1667941163
transform 1 0 37536 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__B1
timestamp 1667941163
transform -1 0 47012 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__A2
timestamp 1667941163
transform 1 0 46828 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__B
timestamp 1667941163
transform -1 0 39468 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__B1
timestamp 1667941163
transform 1 0 39284 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__B
timestamp 1667941163
transform 1 0 34868 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__A1
timestamp 1667941163
transform 1 0 40020 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__A1
timestamp 1667941163
transform -1 0 44160 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__B1
timestamp 1667941163
transform 1 0 51428 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__A1
timestamp 1667941163
transform -1 0 54832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__A1
timestamp 1667941163
transform 1 0 55476 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__B2
timestamp 1667941163
transform -1 0 55384 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__A1
timestamp 1667941163
transform 1 0 52900 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__A1
timestamp 1667941163
transform -1 0 51704 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__B2
timestamp 1667941163
transform 1 0 51980 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A1
timestamp 1667941163
transform 1 0 41952 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__B2
timestamp 1667941163
transform 1 0 44252 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__A1
timestamp 1667941163
transform 1 0 42780 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__B1
timestamp 1667941163
transform 1 0 34132 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__B1
timestamp 1667941163
transform 1 0 34224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__A1
timestamp 1667941163
transform 1 0 52900 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A1
timestamp 1667941163
transform 1 0 52900 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__B2
timestamp 1667941163
transform 1 0 54464 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__A1
timestamp 1667941163
transform -1 0 50508 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__A1
timestamp 1667941163
transform 1 0 52348 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__B2
timestamp 1667941163
transform 1 0 50968 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__A1
timestamp 1667941163
transform 1 0 50324 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__A1
timestamp 1667941163
transform 1 0 50876 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__B1
timestamp 1667941163
transform 1 0 57868 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A1_N
timestamp 1667941163
transform 1 0 52716 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__B2
timestamp 1667941163
transform 1 0 54924 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__A1
timestamp 1667941163
transform 1 0 52072 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__A1
timestamp 1667941163
transform 1 0 54832 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__A1
timestamp 1667941163
transform 1 0 54004 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__B2
timestamp 1667941163
transform 1 0 53452 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__A1
timestamp 1667941163
transform 1 0 55752 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__A1
timestamp 1667941163
transform 1 0 46736 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__A1
timestamp 1667941163
transform 1 0 47840 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__B2
timestamp 1667941163
transform 1 0 50324 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__A1_N
timestamp 1667941163
transform -1 0 58236 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__B2
timestamp 1667941163
transform -1 0 56948 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__A1
timestamp 1667941163
transform 1 0 56764 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__B1
timestamp 1667941163
transform 1 0 56672 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__A1_N
timestamp 1667941163
transform 1 0 56028 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__B2
timestamp 1667941163
transform 1 0 56488 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__A1
timestamp 1667941163
transform 1 0 54280 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__A
timestamp 1667941163
transform -1 0 39284 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__A1
timestamp 1667941163
transform 1 0 50232 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__A1
timestamp 1667941163
transform -1 0 52440 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__B2
timestamp 1667941163
transform 1 0 51704 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__A1
timestamp 1667941163
transform 1 0 49680 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__A1
timestamp 1667941163
transform 1 0 56304 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__B2
timestamp 1667941163
transform 1 0 55752 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__B1
timestamp 1667941163
transform -1 0 58052 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__B1
timestamp 1667941163
transform -1 0 55752 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__A1
timestamp 1667941163
transform -1 0 51520 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__A1
timestamp 1667941163
transform 1 0 52256 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__B2
timestamp 1667941163
transform 1 0 51796 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__A1
timestamp 1667941163
transform 1 0 56028 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__A1
timestamp 1667941163
transform 1 0 56580 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__B2
timestamp 1667941163
transform 1 0 55200 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__A1_N
timestamp 1667941163
transform 1 0 56304 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__B2
timestamp 1667941163
transform -1 0 58236 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__A1
timestamp 1667941163
transform -1 0 57500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__B1_N
timestamp 1667941163
transform -1 0 58236 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__A1_N
timestamp 1667941163
transform 1 0 56488 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__B2
timestamp 1667941163
transform -1 0 55660 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__A1
timestamp 1667941163
transform -1 0 56856 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__A1
timestamp 1667941163
transform -1 0 47932 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__A1
timestamp 1667941163
transform 1 0 45632 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__B2
timestamp 1667941163
transform 1 0 49680 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__A
timestamp 1667941163
transform 1 0 43700 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__A1
timestamp 1667941163
transform 1 0 55752 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__A1
timestamp 1667941163
transform 1 0 54648 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__B2
timestamp 1667941163
transform 1 0 53176 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__B1
timestamp 1667941163
transform -1 0 58236 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__A1
timestamp 1667941163
transform -1 0 51244 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__A1
timestamp 1667941163
transform 1 0 51980 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__B2
timestamp 1667941163
transform 1 0 52532 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__A1
timestamp 1667941163
transform 1 0 55292 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__A1
timestamp 1667941163
transform 1 0 57316 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__B2
timestamp 1667941163
transform 1 0 56488 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__A1_N
timestamp 1667941163
transform 1 0 56580 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__B2
timestamp 1667941163
transform 1 0 54188 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__A1
timestamp 1667941163
transform -1 0 53636 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__A1
timestamp 1667941163
transform 1 0 49220 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__A1
timestamp 1667941163
transform -1 0 49312 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__B2
timestamp 1667941163
transform 1 0 49404 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__A1
timestamp 1667941163
transform 1 0 54004 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__A1
timestamp 1667941163
transform 1 0 55016 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__B2
timestamp 1667941163
transform 1 0 54464 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__A1_N
timestamp 1667941163
transform -1 0 58236 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__B2
timestamp 1667941163
transform -1 0 58236 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__A1
timestamp 1667941163
transform -1 0 56212 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__A1
timestamp 1667941163
transform -1 0 58236 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__A1
timestamp 1667941163
transform 1 0 57224 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__B2
timestamp 1667941163
transform 1 0 51428 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__A
timestamp 1667941163
transform 1 0 49680 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1504__A1
timestamp 1667941163
transform 1 0 49680 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1504__B2
timestamp 1667941163
transform 1 0 49772 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__B2
timestamp 1667941163
transform 1 0 50784 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1509__A
timestamp 1667941163
transform 1 0 47104 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1511__A1_N
timestamp 1667941163
transform -1 0 55660 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1511__B2
timestamp 1667941163
transform -1 0 58144 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__A1
timestamp 1667941163
transform -1 0 56212 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__A1
timestamp 1667941163
transform -1 0 47932 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__A1
timestamp 1667941163
transform 1 0 49772 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__B2
timestamp 1667941163
transform 1 0 48576 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1520__A1
timestamp 1667941163
transform 1 0 52256 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__A1
timestamp 1667941163
transform 1 0 56120 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__B2
timestamp 1667941163
transform 1 0 54556 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1524__A1
timestamp 1667941163
transform 1 0 52164 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1524__B2
timestamp 1667941163
transform 1 0 51336 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1525__A1
timestamp 1667941163
transform 1 0 52716 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1528__A1_N
timestamp 1667941163
transform -1 0 55844 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1528__B2
timestamp 1667941163
transform -1 0 55292 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1529__A1
timestamp 1667941163
transform -1 0 54740 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1534__A1_N
timestamp 1667941163
transform 1 0 56304 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1534__B2
timestamp 1667941163
transform -1 0 53728 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__A1
timestamp 1667941163
transform 1 0 52900 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1539__A1_N
timestamp 1667941163
transform -1 0 58420 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1539__B2
timestamp 1667941163
transform -1 0 57224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1540__A1
timestamp 1667941163
transform -1 0 56396 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1545__S
timestamp 1667941163
transform 1 0 54372 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1550__A1_N
timestamp 1667941163
transform 1 0 51704 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1555__A1
timestamp 1667941163
transform 1 0 51152 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1556__A1
timestamp 1667941163
transform 1 0 50968 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1556__B2
timestamp 1667941163
transform 1 0 53268 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1559__B1_N
timestamp 1667941163
transform 1 0 51520 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1560__A1
timestamp 1667941163
transform 1 0 50416 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1563__B1
timestamp 1667941163
transform 1 0 47748 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1565__A1
timestamp 1667941163
transform 1 0 53360 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1575__S
timestamp 1667941163
transform 1 0 47104 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1578__A1
timestamp 1667941163
transform -1 0 51152 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1578__S0
timestamp 1667941163
transform -1 0 47932 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1579__S
timestamp 1667941163
transform 1 0 51612 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1580__A1
timestamp 1667941163
transform -1 0 52164 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1583__A1
timestamp 1667941163
transform 1 0 50324 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1586__A1
timestamp 1667941163
transform -1 0 52164 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1600__CLK
timestamp 1667941163
transform -1 0 40572 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1602__CLK
timestamp 1667941163
transform 1 0 42596 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1604__CLK
timestamp 1667941163
transform -1 0 38916 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1614__CLK
timestamp 1667941163
transform -1 0 44620 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1615__CLK
timestamp 1667941163
transform 1 0 34408 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1624__CLK
timestamp 1667941163
transform 1 0 46000 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1626__CLK
timestamp 1667941163
transform 1 0 46552 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1633__CLK
timestamp 1667941163
transform 1 0 34224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1637__CLK
timestamp 1667941163
transform 1 0 35420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1638__CLK
timestamp 1667941163
transform 1 0 37812 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout8_A
timestamp 1667941163
transform 1 0 29348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout9_A
timestamp 1667941163
transform 1 0 27508 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout10_A
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout11_A
timestamp 1667941163
transform 1 0 46828 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout12_A
timestamp 1667941163
transform -1 0 47932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout13_A
timestamp 1667941163
transform -1 0 44436 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform -1 0 58420 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1667941163
transform -1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1667941163
transform -1 0 1748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1667941163
transform -1 0 3128 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1667941163
transform -1 0 58420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output7_A
timestamp 1667941163
transform -1 0 2484 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9 OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1667941163
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1667941163
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1667941163
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1667941163
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1667941163
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1667941163
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1667941163
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1667941163
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1667941163
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1667941163
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1667941163
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1667941163
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1667941163
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1667941163
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_293 OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28060 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_301
timestamp 1667941163
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1667941163
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_315
timestamp 1667941163
transform 1 0 30084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1667941163
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1667941163
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1667941163
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1667941163
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1667941163
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1667941163
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1667941163
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1667941163
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1667941163
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1667941163
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1667941163
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1667941163
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1667941163
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1667941163
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1667941163
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1667941163
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1667941163
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1667941163
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1667941163
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1667941163
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1667941163
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1667941163
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1667941163
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1667941163
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1667941163
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_617
timestamp 1667941163
transform 1 0 57868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_623
timestamp 1667941163
transform 1 0 58420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7
timestamp 1667941163
transform 1 0 1748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1667941163
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1667941163
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_43
timestamp 1667941163
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1667941163
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1667941163
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1667941163
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1667941163
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1667941163
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1667941163
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1667941163
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1667941163
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1667941163
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1667941163
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1667941163
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1667941163
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1667941163
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1667941163
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1667941163
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1667941163
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1667941163
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1667941163
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1667941163
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1667941163
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1667941163
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1667941163
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1667941163
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1667941163
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1667941163
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1667941163
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1667941163
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1667941163
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1667941163
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_617 OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 57868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_623
timestamp 1667941163
transform 1 0 58420 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1667941163
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1667941163
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1667941163
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1667941163
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1667941163
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1667941163
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1667941163
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1667941163
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1667941163
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1667941163
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1667941163
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1667941163
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1667941163
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1667941163
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1667941163
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1667941163
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1667941163
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1667941163
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1667941163
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1667941163
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1667941163
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1667941163
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1667941163
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1667941163
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1667941163
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1667941163
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1667941163
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1667941163
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1667941163
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1667941163
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1667941163
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1667941163
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1667941163
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1667941163
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1667941163
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1667941163
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1667941163
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1667941163
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1667941163
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1667941163
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1667941163
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1667941163
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1667941163
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1667941163
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1667941163
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1667941163
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_617
timestamp 1667941163
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1667941163
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1667941163
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1667941163
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1667941163
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1667941163
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1667941163
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1667941163
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1667941163
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1667941163
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1667941163
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1667941163
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1667941163
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1667941163
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1667941163
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1667941163
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1667941163
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1667941163
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1667941163
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1667941163
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1667941163
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1667941163
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1667941163
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1667941163
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1667941163
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1667941163
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1667941163
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1667941163
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1667941163
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1667941163
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1667941163
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1667941163
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1667941163
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1667941163
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1667941163
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1667941163
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1667941163
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1667941163
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1667941163
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1667941163
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1667941163
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1667941163
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1667941163
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1667941163
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1667941163
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1667941163
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1667941163
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1667941163
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1667941163
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1667941163
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1667941163
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1667941163
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1667941163
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1667941163
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1667941163
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1667941163
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1667941163
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1667941163
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1667941163
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1667941163
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1667941163
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1667941163
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1667941163
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1667941163
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1667941163
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1667941163
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1667941163
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1667941163
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1667941163
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1667941163
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1667941163
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1667941163
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1667941163
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1667941163
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1667941163
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1667941163
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1667941163
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1667941163
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1667941163
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1667941163
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1667941163
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1667941163
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1667941163
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1667941163
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1667941163
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1667941163
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1667941163
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1667941163
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1667941163
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1667941163
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1667941163
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1667941163
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1667941163
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1667941163
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1667941163
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1667941163
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1667941163
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1667941163
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1667941163
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1667941163
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1667941163
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1667941163
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1667941163
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1667941163
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1667941163
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1667941163
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1667941163
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1667941163
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1667941163
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1667941163
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1667941163
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1667941163
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1667941163
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1667941163
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1667941163
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1667941163
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1667941163
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1667941163
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1667941163
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1667941163
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1667941163
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1667941163
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1667941163
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1667941163
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1667941163
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1667941163
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1667941163
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1667941163
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1667941163
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1667941163
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1667941163
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1667941163
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1667941163
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1667941163
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1667941163
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1667941163
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1667941163
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1667941163
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1667941163
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1667941163
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1667941163
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1667941163
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1667941163
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1667941163
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1667941163
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1667941163
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1667941163
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1667941163
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1667941163
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1667941163
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1667941163
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1667941163
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1667941163
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1667941163
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1667941163
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1667941163
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1667941163
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1667941163
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1667941163
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1667941163
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1667941163
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1667941163
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1667941163
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1667941163
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1667941163
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1667941163
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1667941163
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1667941163
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1667941163
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1667941163
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1667941163
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1667941163
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1667941163
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1667941163
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1667941163
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1667941163
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1667941163
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1667941163
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1667941163
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1667941163
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1667941163
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1667941163
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1667941163
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1667941163
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1667941163
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1667941163
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1667941163
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1667941163
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1667941163
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1667941163
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1667941163
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1667941163
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1667941163
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1667941163
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1667941163
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1667941163
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1667941163
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1667941163
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1667941163
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1667941163
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1667941163
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1667941163
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1667941163
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1667941163
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1667941163
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1667941163
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1667941163
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1667941163
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1667941163
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1667941163
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1667941163
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1667941163
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1667941163
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1667941163
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1667941163
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1667941163
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1667941163
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1667941163
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1667941163
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1667941163
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1667941163
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1667941163
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1667941163
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1667941163
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1667941163
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1667941163
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1667941163
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1667941163
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1667941163
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1667941163
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1667941163
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1667941163
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1667941163
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1667941163
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1667941163
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1667941163
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1667941163
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1667941163
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1667941163
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1667941163
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1667941163
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1667941163
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1667941163
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1667941163
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1667941163
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1667941163
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1667941163
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1667941163
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1667941163
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1667941163
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1667941163
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1667941163
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1667941163
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1667941163
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1667941163
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1667941163
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1667941163
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1667941163
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1667941163
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1667941163
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1667941163
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1667941163
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1667941163
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1667941163
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1667941163
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1667941163
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1667941163
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1667941163
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1667941163
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1667941163
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1667941163
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1667941163
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1667941163
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1667941163
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1667941163
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1667941163
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1667941163
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1667941163
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1667941163
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1667941163
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1667941163
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1667941163
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1667941163
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1667941163
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1667941163
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1667941163
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1667941163
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1667941163
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1667941163
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1667941163
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1667941163
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1667941163
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1667941163
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1667941163
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1667941163
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1667941163
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1667941163
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1667941163
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1667941163
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1667941163
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1667941163
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1667941163
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1667941163
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1667941163
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1667941163
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1667941163
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1667941163
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1667941163
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1667941163
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1667941163
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1667941163
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1667941163
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1667941163
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1667941163
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1667941163
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1667941163
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1667941163
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1667941163
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1667941163
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1667941163
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1667941163
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1667941163
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1667941163
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1667941163
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1667941163
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1667941163
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1667941163
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1667941163
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1667941163
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1667941163
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1667941163
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1667941163
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1667941163
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1667941163
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1667941163
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1667941163
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1667941163
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1667941163
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1667941163
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1667941163
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1667941163
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1667941163
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1667941163
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1667941163
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1667941163
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1667941163
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1667941163
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1667941163
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1667941163
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1667941163
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1667941163
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1667941163
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1667941163
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1667941163
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1667941163
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1667941163
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1667941163
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1667941163
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1667941163
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1667941163
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1667941163
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1667941163
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1667941163
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1667941163
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1667941163
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1667941163
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1667941163
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1667941163
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1667941163
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1667941163
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1667941163
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1667941163
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1667941163
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1667941163
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1667941163
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1667941163
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1667941163
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1667941163
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1667941163
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1667941163
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1667941163
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1667941163
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1667941163
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1667941163
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1667941163
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1667941163
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1667941163
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1667941163
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1667941163
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1667941163
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1667941163
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1667941163
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1667941163
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1667941163
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1667941163
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1667941163
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1667941163
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1667941163
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1667941163
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1667941163
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1667941163
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1667941163
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1667941163
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1667941163
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1667941163
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1667941163
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1667941163
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1667941163
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1667941163
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1667941163
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1667941163
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1667941163
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1667941163
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1667941163
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1667941163
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1667941163
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1667941163
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1667941163
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1667941163
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1667941163
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1667941163
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1667941163
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1667941163
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1667941163
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1667941163
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1667941163
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1667941163
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1667941163
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1667941163
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1667941163
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1667941163
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1667941163
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1667941163
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1667941163
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1667941163
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1667941163
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1667941163
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1667941163
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1667941163
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1667941163
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1667941163
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1667941163
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1667941163
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1667941163
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1667941163
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1667941163
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1667941163
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1667941163
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1667941163
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1667941163
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1667941163
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1667941163
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1667941163
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1667941163
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1667941163
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1667941163
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1667941163
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1667941163
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1667941163
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1667941163
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1667941163
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1667941163
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1667941163
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1667941163
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1667941163
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1667941163
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1667941163
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1667941163
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1667941163
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1667941163
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1667941163
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1667941163
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1667941163
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1667941163
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1667941163
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1667941163
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1667941163
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1667941163
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1667941163
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1667941163
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1667941163
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1667941163
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1667941163
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1667941163
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1667941163
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1667941163
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1667941163
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1667941163
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1667941163
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1667941163
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1667941163
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1667941163
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1667941163
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1667941163
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1667941163
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1667941163
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1667941163
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1667941163
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1667941163
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1667941163
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1667941163
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1667941163
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1667941163
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1667941163
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1667941163
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1667941163
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1667941163
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1667941163
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1667941163
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1667941163
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1667941163
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1667941163
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1667941163
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1667941163
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1667941163
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1667941163
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1667941163
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1667941163
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1667941163
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1667941163
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1667941163
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1667941163
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1667941163
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1667941163
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1667941163
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1667941163
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1667941163
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1667941163
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1667941163
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1667941163
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1667941163
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1667941163
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1667941163
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1667941163
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1667941163
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1667941163
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1667941163
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1667941163
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1667941163
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1667941163
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1667941163
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1667941163
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1667941163
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1667941163
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1667941163
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1667941163
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1667941163
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1667941163
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1667941163
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1667941163
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1667941163
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1667941163
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1667941163
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1667941163
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1667941163
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1667941163
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1667941163
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1667941163
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1667941163
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1667941163
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1667941163
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1667941163
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1667941163
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1667941163
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1667941163
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1667941163
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1667941163
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1667941163
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1667941163
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1667941163
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1667941163
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1667941163
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1667941163
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1667941163
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1667941163
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1667941163
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1667941163
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1667941163
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1667941163
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1667941163
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1667941163
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1667941163
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1667941163
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1667941163
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1667941163
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1667941163
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1667941163
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1667941163
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1667941163
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1667941163
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1667941163
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1667941163
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1667941163
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1667941163
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1667941163
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1667941163
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1667941163
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1667941163
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1667941163
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1667941163
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1667941163
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1667941163
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1667941163
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1667941163
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1667941163
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1667941163
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1667941163
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1667941163
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1667941163
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1667941163
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1667941163
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1667941163
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1667941163
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1667941163
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1667941163
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1667941163
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1667941163
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1667941163
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1667941163
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1667941163
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1667941163
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1667941163
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1667941163
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1667941163
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1667941163
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1667941163
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1667941163
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1667941163
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1667941163
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1667941163
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1667941163
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1667941163
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1667941163
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1667941163
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1667941163
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1667941163
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1667941163
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1667941163
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1667941163
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1667941163
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1667941163
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1667941163
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1667941163
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1667941163
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1667941163
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1667941163
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1667941163
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1667941163
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1667941163
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1667941163
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1667941163
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1667941163
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1667941163
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1667941163
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1667941163
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1667941163
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1667941163
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1667941163
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1667941163
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1667941163
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1667941163
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1667941163
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1667941163
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1667941163
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1667941163
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1667941163
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1667941163
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1667941163
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1667941163
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1667941163
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1667941163
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1667941163
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1667941163
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1667941163
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1667941163
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1667941163
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1667941163
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1667941163
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1667941163
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1667941163
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1667941163
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1667941163
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1667941163
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1667941163
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1667941163
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1667941163
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1667941163
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1667941163
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1667941163
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1667941163
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1667941163
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1667941163
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1667941163
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1667941163
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1667941163
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1667941163
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1667941163
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1667941163
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1667941163
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1667941163
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1667941163
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1667941163
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1667941163
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1667941163
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1667941163
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1667941163
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1667941163
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1667941163
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1667941163
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1667941163
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1667941163
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1667941163
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1667941163
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1667941163
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1667941163
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1667941163
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1667941163
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1667941163
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1667941163
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1667941163
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1667941163
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1667941163
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1667941163
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1667941163
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1667941163
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1667941163
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1667941163
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1667941163
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1667941163
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1667941163
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1667941163
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1667941163
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1667941163
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1667941163
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1667941163
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1667941163
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1667941163
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1667941163
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1667941163
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1667941163
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1667941163
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1667941163
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1667941163
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1667941163
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1667941163
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1667941163
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1667941163
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1667941163
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1667941163
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1667941163
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1667941163
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1667941163
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1667941163
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1667941163
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1667941163
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1667941163
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1667941163
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1667941163
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1667941163
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1667941163
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1667941163
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1667941163
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1667941163
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1667941163
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1667941163
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1667941163
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1667941163
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1667941163
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1667941163
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1667941163
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1667941163
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1667941163
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1667941163
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1667941163
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1667941163
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1667941163
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1667941163
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1667941163
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1667941163
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1667941163
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1667941163
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1667941163
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1667941163
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1667941163
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1667941163
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1667941163
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1667941163
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1667941163
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1667941163
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1667941163
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1667941163
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1667941163
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1667941163
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1667941163
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1667941163
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1667941163
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1667941163
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1667941163
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1667941163
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1667941163
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1667941163
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1667941163
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1667941163
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1667941163
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1667941163
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1667941163
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1667941163
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1667941163
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1667941163
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1667941163
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1667941163
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1667941163
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1667941163
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1667941163
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1667941163
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1667941163
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1667941163
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1667941163
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1667941163
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1667941163
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1667941163
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1667941163
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1667941163
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1667941163
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1667941163
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1667941163
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1667941163
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_489
timestamp 1667941163
transform 1 0 46092 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_517
timestamp 1667941163
transform 1 0 48668 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_529
timestamp 1667941163
transform 1 0 49772 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1667941163
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1667941163
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1667941163
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1667941163
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1667941163
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1667941163
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1667941163
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1667941163
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1667941163
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1667941163
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1667941163
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1667941163
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1667941163
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1667941163
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1667941163
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_398
timestamp 1667941163
transform 1 0 37720 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_416
timestamp 1667941163
transform 1 0 39376 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_428
timestamp 1667941163
transform 1 0 40480 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_440
timestamp 1667941163
transform 1 0 41584 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1667941163
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1667941163
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1667941163
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1667941163
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1667941163
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1667941163
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_505
timestamp 1667941163
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_509
timestamp 1667941163
transform 1 0 47932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_521
timestamp 1667941163
transform 1 0 49036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_533
timestamp 1667941163
transform 1 0 50140 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_545
timestamp 1667941163
transform 1 0 51244 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_557
timestamp 1667941163
transform 1 0 52348 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1667941163
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1667941163
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1667941163
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1667941163
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1667941163
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1667941163
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_617
timestamp 1667941163
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1667941163
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_375
timestamp 1667941163
transform 1 0 35604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_402
timestamp 1667941163
transform 1 0 38088 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_409
timestamp 1667941163
transform 1 0 38732 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1667941163
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1667941163
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1667941163
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1667941163
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1667941163
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1667941163
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1667941163
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1667941163
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1667941163
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_504
timestamp 1667941163
transform 1 0 47472 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_511
timestamp 1667941163
transform 1 0 48116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_518
timestamp 1667941163
transform 1 0 48760 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1667941163
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1667941163
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1667941163
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1667941163
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1667941163
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1667941163
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1667941163
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1667941163
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1667941163
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1667941163
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1667941163
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1667941163
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1667941163
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1667941163
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1667941163
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1667941163
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_379
timestamp 1667941163
transform 1 0 35972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_383
timestamp 1667941163
transform 1 0 36340 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1667941163
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_398
timestamp 1667941163
transform 1 0 37720 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_422
timestamp 1667941163
transform 1 0 39928 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_433
timestamp 1667941163
transform 1 0 40940 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_439
timestamp 1667941163
transform 1 0 41492 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1667941163
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1667941163
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_461
timestamp 1667941163
transform 1 0 43516 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_467
timestamp 1667941163
transform 1 0 44068 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_491
timestamp 1667941163
transform 1 0 46276 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_498
timestamp 1667941163
transform 1 0 46920 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_505
timestamp 1667941163
transform 1 0 47564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_509
timestamp 1667941163
transform 1 0 47932 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_530
timestamp 1667941163
transform 1 0 49864 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_538
timestamp 1667941163
transform 1 0 50600 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_545
timestamp 1667941163
transform 1 0 51244 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_551
timestamp 1667941163
transform 1 0 51796 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1667941163
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1667941163
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1667941163
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1667941163
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1667941163
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1667941163
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1667941163
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_617
timestamp 1667941163
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1667941163
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1667941163
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1667941163
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1667941163
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_381
timestamp 1667941163
transform 1 0 36156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_395
timestamp 1667941163
transform 1 0 37444 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_409
timestamp 1667941163
transform 1 0 38732 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_417
timestamp 1667941163
transform 1 0 39468 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1667941163
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_446
timestamp 1667941163
transform 1 0 42136 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_456
timestamp 1667941163
transform 1 0 43056 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_467
timestamp 1667941163
transform 1 0 44068 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_474
timestamp 1667941163
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_477
timestamp 1667941163
transform 1 0 44988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_482
timestamp 1667941163
transform 1 0 45448 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_510
timestamp 1667941163
transform 1 0 48024 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1667941163
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1667941163
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_533
timestamp 1667941163
transform 1 0 50140 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_555
timestamp 1667941163
transform 1 0 52164 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_567
timestamp 1667941163
transform 1 0 53268 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_579
timestamp 1667941163
transform 1 0 54372 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1667941163
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1667941163
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1667941163
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1667941163
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1667941163
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1667941163
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_357
timestamp 1667941163
transform 1 0 33948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_362
timestamp 1667941163
transform 1 0 34408 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_387
timestamp 1667941163
transform 1 0 36708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_403
timestamp 1667941163
transform 1 0 38180 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_411
timestamp 1667941163
transform 1 0 38916 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_421
timestamp 1667941163
transform 1 0 39836 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_446
timestamp 1667941163
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_449
timestamp 1667941163
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_454
timestamp 1667941163
transform 1 0 42872 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_461
timestamp 1667941163
transform 1 0 43516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_465
timestamp 1667941163
transform 1 0 43884 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_489
timestamp 1667941163
transform 1 0 46092 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_496
timestamp 1667941163
transform 1 0 46736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_502
timestamp 1667941163
transform 1 0 47288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_505
timestamp 1667941163
transform 1 0 47564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_517
timestamp 1667941163
transform 1 0 48668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_524
timestamp 1667941163
transform 1 0 49312 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_528
timestamp 1667941163
transform 1 0 49680 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_552
timestamp 1667941163
transform 1 0 51888 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1667941163
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1667941163
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1667941163
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1667941163
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1667941163
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1667941163
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1667941163
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1667941163
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_372
timestamp 1667941163
transform 1 0 35328 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_379
timestamp 1667941163
transform 1 0 35972 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_385
timestamp 1667941163
transform 1 0 36524 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_395
timestamp 1667941163
transform 1 0 37444 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_406
timestamp 1667941163
transform 1 0 38456 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1667941163
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1667941163
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_444
timestamp 1667941163
transform 1 0 41952 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_450
timestamp 1667941163
transform 1 0 42504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_455
timestamp 1667941163
transform 1 0 42964 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_462
timestamp 1667941163
transform 1 0 43608 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_468
timestamp 1667941163
transform 1 0 44160 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_474
timestamp 1667941163
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1667941163
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_482
timestamp 1667941163
transform 1 0 45448 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_490
timestamp 1667941163
transform 1 0 46184 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_495
timestamp 1667941163
transform 1 0 46644 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_523
timestamp 1667941163
transform 1 0 49220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_529
timestamp 1667941163
transform 1 0 49772 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_533
timestamp 1667941163
transform 1 0 50140 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_542
timestamp 1667941163
transform 1 0 50968 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_549
timestamp 1667941163
transform 1 0 51612 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_561
timestamp 1667941163
transform 1 0 52716 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_573
timestamp 1667941163
transform 1 0 53820 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_585
timestamp 1667941163
transform 1 0 54924 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1667941163
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1667941163
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1667941163
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1667941163
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1667941163
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1667941163
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1667941163
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1667941163
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_384
timestamp 1667941163
transform 1 0 36432 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_403
timestamp 1667941163
transform 1 0 38180 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_409
timestamp 1667941163
transform 1 0 38732 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_415
timestamp 1667941163
transform 1 0 39284 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_424
timestamp 1667941163
transform 1 0 40112 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_435
timestamp 1667941163
transform 1 0 41124 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_443
timestamp 1667941163
transform 1 0 41860 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1667941163
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_449
timestamp 1667941163
transform 1 0 42412 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_455
timestamp 1667941163
transform 1 0 42964 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_463
timestamp 1667941163
transform 1 0 43700 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_487
timestamp 1667941163
transform 1 0 45908 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_498
timestamp 1667941163
transform 1 0 46920 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_505
timestamp 1667941163
transform 1 0 47564 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_509
timestamp 1667941163
transform 1 0 47932 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_517
timestamp 1667941163
transform 1 0 48668 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_538
timestamp 1667941163
transform 1 0 50600 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_549
timestamp 1667941163
transform 1 0 51612 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_557
timestamp 1667941163
transform 1 0 52348 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1667941163
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1667941163
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1667941163
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1667941163
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1667941163
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1667941163
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1667941163
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1667941163
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1667941163
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1667941163
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1667941163
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1667941163
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_369
timestamp 1667941163
transform 1 0 35052 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_376
timestamp 1667941163
transform 1 0 35696 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_387
timestamp 1667941163
transform 1 0 36708 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_397
timestamp 1667941163
transform 1 0 37628 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_407
timestamp 1667941163
transform 1 0 38548 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_416
timestamp 1667941163
transform 1 0 39376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_421
timestamp 1667941163
transform 1 0 39836 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_431
timestamp 1667941163
transform 1 0 40756 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_456
timestamp 1667941163
transform 1 0 43056 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_462
timestamp 1667941163
transform 1 0 43608 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_468
timestamp 1667941163
transform 1 0 44160 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_474
timestamp 1667941163
transform 1 0 44712 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_477
timestamp 1667941163
transform 1 0 44988 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_482
timestamp 1667941163
transform 1 0 45448 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_490
timestamp 1667941163
transform 1 0 46184 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_494
timestamp 1667941163
transform 1 0 46552 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_505
timestamp 1667941163
transform 1 0 47564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_514
timestamp 1667941163
transform 1 0 48392 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_518
timestamp 1667941163
transform 1 0 48760 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_523
timestamp 1667941163
transform 1 0 49220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_529
timestamp 1667941163
transform 1 0 49772 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_533
timestamp 1667941163
transform 1 0 50140 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_537
timestamp 1667941163
transform 1 0 50508 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_541
timestamp 1667941163
transform 1 0 50876 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_561
timestamp 1667941163
transform 1 0 52716 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_573
timestamp 1667941163
transform 1 0 53820 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1667941163
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1667941163
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1667941163
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1667941163
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1667941163
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1667941163
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_364
timestamp 1667941163
transform 1 0 34592 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_371
timestamp 1667941163
transform 1 0 35236 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_386
timestamp 1667941163
transform 1 0 36616 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_401
timestamp 1667941163
transform 1 0 37996 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_408
timestamp 1667941163
transform 1 0 38640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_420
timestamp 1667941163
transform 1 0 39744 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_446
timestamp 1667941163
transform 1 0 42136 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_449
timestamp 1667941163
transform 1 0 42412 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_457
timestamp 1667941163
transform 1 0 43148 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_464
timestamp 1667941163
transform 1 0 43792 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_468
timestamp 1667941163
transform 1 0 44160 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_472
timestamp 1667941163
transform 1 0 44528 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_478
timestamp 1667941163
transform 1 0 45080 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_486
timestamp 1667941163
transform 1 0 45816 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_493
timestamp 1667941163
transform 1 0 46460 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_499
timestamp 1667941163
transform 1 0 47012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1667941163
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_505
timestamp 1667941163
transform 1 0 47564 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_515
timestamp 1667941163
transform 1 0 48484 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_524
timestamp 1667941163
transform 1 0 49312 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_531
timestamp 1667941163
transform 1 0 49956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_537
timestamp 1667941163
transform 1 0 50508 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_543
timestamp 1667941163
transform 1 0 51060 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_549
timestamp 1667941163
transform 1 0 51612 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_555
timestamp 1667941163
transform 1 0 52164 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1667941163
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_561
timestamp 1667941163
transform 1 0 52716 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_569
timestamp 1667941163
transform 1 0 53452 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_572
timestamp 1667941163
transform 1 0 53728 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_580
timestamp 1667941163
transform 1 0 54464 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_583
timestamp 1667941163
transform 1 0 54740 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_589
timestamp 1667941163
transform 1 0 55292 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_595
timestamp 1667941163
transform 1 0 55844 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_601
timestamp 1667941163
transform 1 0 56396 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_613
timestamp 1667941163
transform 1 0 57500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1667941163
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1667941163
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1667941163
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1667941163
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1667941163
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1667941163
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_347
timestamp 1667941163
transform 1 0 33028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1667941163
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_387
timestamp 1667941163
transform 1 0 36708 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_407
timestamp 1667941163
transform 1 0 38548 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_418
timestamp 1667941163
transform 1 0 39560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_421
timestamp 1667941163
transform 1 0 39836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_430
timestamp 1667941163
transform 1 0 40664 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_434
timestamp 1667941163
transform 1 0 41032 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_444
timestamp 1667941163
transform 1 0 41952 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1667941163
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1667941163
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_477
timestamp 1667941163
transform 1 0 44988 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_482
timestamp 1667941163
transform 1 0 45448 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_495
timestamp 1667941163
transform 1 0 46644 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_502
timestamp 1667941163
transform 1 0 47288 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_506
timestamp 1667941163
transform 1 0 47656 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_511
timestamp 1667941163
transform 1 0 48116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_518
timestamp 1667941163
transform 1 0 48760 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_530
timestamp 1667941163
transform 1 0 49864 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_533
timestamp 1667941163
transform 1 0 50140 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_538
timestamp 1667941163
transform 1 0 50600 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_559
timestamp 1667941163
transform 1 0 52532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_565
timestamp 1667941163
transform 1 0 53084 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_571
timestamp 1667941163
transform 1 0 53636 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_583
timestamp 1667941163
transform 1 0 54740 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1667941163
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_589
timestamp 1667941163
transform 1 0 55292 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_593
timestamp 1667941163
transform 1 0 55660 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_599
timestamp 1667941163
transform 1 0 56212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_603
timestamp 1667941163
transform 1 0 56580 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_606
timestamp 1667941163
transform 1 0 56856 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_612
timestamp 1667941163
transform 1 0 57408 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_624
timestamp 1667941163
transform 1 0 58512 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_345
timestamp 1667941163
transform 1 0 32844 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_371
timestamp 1667941163
transform 1 0 35236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_384
timestamp 1667941163
transform 1 0 36432 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_390
timestamp 1667941163
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_401
timestamp 1667941163
transform 1 0 37996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_413
timestamp 1667941163
transform 1 0 39100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_420
timestamp 1667941163
transform 1 0 39744 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_446
timestamp 1667941163
transform 1 0 42136 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_449
timestamp 1667941163
transform 1 0 42412 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_457
timestamp 1667941163
transform 1 0 43148 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_461
timestamp 1667941163
transform 1 0 43516 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_468
timestamp 1667941163
transform 1 0 44160 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_478
timestamp 1667941163
transform 1 0 45080 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_484
timestamp 1667941163
transform 1 0 45632 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_495
timestamp 1667941163
transform 1 0 46644 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_502
timestamp 1667941163
transform 1 0 47288 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_505
timestamp 1667941163
transform 1 0 47564 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_510
timestamp 1667941163
transform 1 0 48024 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_523
timestamp 1667941163
transform 1 0 49220 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_531
timestamp 1667941163
transform 1 0 49956 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_540
timestamp 1667941163
transform 1 0 50784 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_551
timestamp 1667941163
transform 1 0 51796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_557
timestamp 1667941163
transform 1 0 52348 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_561
timestamp 1667941163
transform 1 0 52716 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_565
timestamp 1667941163
transform 1 0 53084 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_573
timestamp 1667941163
transform 1 0 53820 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_579
timestamp 1667941163
transform 1 0 54372 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_590
timestamp 1667941163
transform 1 0 55384 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_598
timestamp 1667941163
transform 1 0 56120 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_604
timestamp 1667941163
transform 1 0 56672 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_610
timestamp 1667941163
transform 1 0 57224 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_617
timestamp 1667941163
transform 1 0 57868 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_621
timestamp 1667941163
transform 1 0 58236 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_341
timestamp 1667941163
transform 1 0 32476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_356
timestamp 1667941163
transform 1 0 33856 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1667941163
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_380
timestamp 1667941163
transform 1 0 36064 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_386
timestamp 1667941163
transform 1 0 36616 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_394
timestamp 1667941163
transform 1 0 37352 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_402
timestamp 1667941163
transform 1 0 38088 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_410
timestamp 1667941163
transform 1 0 38824 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_418
timestamp 1667941163
transform 1 0 39560 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_421
timestamp 1667941163
transform 1 0 39836 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_428
timestamp 1667941163
transform 1 0 40480 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_436
timestamp 1667941163
transform 1 0 41216 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_440
timestamp 1667941163
transform 1 0 41584 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_461
timestamp 1667941163
transform 1 0 43516 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_468
timestamp 1667941163
transform 1 0 44160 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_474
timestamp 1667941163
transform 1 0 44712 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_477
timestamp 1667941163
transform 1 0 44988 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_485
timestamp 1667941163
transform 1 0 45724 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_495
timestamp 1667941163
transform 1 0 46644 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_503
timestamp 1667941163
transform 1 0 47380 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_509
timestamp 1667941163
transform 1 0 47932 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_518
timestamp 1667941163
transform 1 0 48760 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_527
timestamp 1667941163
transform 1 0 49588 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1667941163
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_533
timestamp 1667941163
transform 1 0 50140 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_540
timestamp 1667941163
transform 1 0 50784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_553
timestamp 1667941163
transform 1 0 51980 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_566
timestamp 1667941163
transform 1 0 53176 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_579
timestamp 1667941163
transform 1 0 54372 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_586
timestamp 1667941163
transform 1 0 55016 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_589
timestamp 1667941163
transform 1 0 55292 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_596
timestamp 1667941163
transform 1 0 55936 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_602
timestamp 1667941163
transform 1 0 56488 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_617
timestamp 1667941163
transform 1 0 57868 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_623
timestamp 1667941163
transform 1 0 58420 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_334
timestamp 1667941163
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_362
timestamp 1667941163
transform 1 0 34408 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_386
timestamp 1667941163
transform 1 0 36616 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_399
timestamp 1667941163
transform 1 0 37812 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_403
timestamp 1667941163
transform 1 0 38180 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_411
timestamp 1667941163
transform 1 0 38916 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_419
timestamp 1667941163
transform 1 0 39652 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_425
timestamp 1667941163
transform 1 0 40204 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_433
timestamp 1667941163
transform 1 0 40940 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_443
timestamp 1667941163
transform 1 0 41860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1667941163
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_449
timestamp 1667941163
transform 1 0 42412 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_454
timestamp 1667941163
transform 1 0 42872 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_460
timestamp 1667941163
transform 1 0 43424 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_464
timestamp 1667941163
transform 1 0 43792 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_473
timestamp 1667941163
transform 1 0 44620 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_486
timestamp 1667941163
transform 1 0 45816 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_498
timestamp 1667941163
transform 1 0 46920 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_505
timestamp 1667941163
transform 1 0 47564 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_510
timestamp 1667941163
transform 1 0 48024 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_523
timestamp 1667941163
transform 1 0 49220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_529
timestamp 1667941163
transform 1 0 49772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_537
timestamp 1667941163
transform 1 0 50508 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_549
timestamp 1667941163
transform 1 0 51612 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_555
timestamp 1667941163
transform 1 0 52164 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1667941163
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_561
timestamp 1667941163
transform 1 0 52716 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_572
timestamp 1667941163
transform 1 0 53728 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_580
timestamp 1667941163
transform 1 0 54464 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_588
timestamp 1667941163
transform 1 0 55200 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_596
timestamp 1667941163
transform 1 0 55936 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_602
timestamp 1667941163
transform 1 0 56488 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_606
timestamp 1667941163
transform 1 0 56856 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_614
timestamp 1667941163
transform 1 0 57592 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_617
timestamp 1667941163
transform 1 0 57868 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_623
timestamp 1667941163
transform 1 0 58420 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1667941163
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1667941163
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1667941163
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1667941163
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_343
timestamp 1667941163
transform 1 0 32660 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_350
timestamp 1667941163
transform 1 0 33304 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_356
timestamp 1667941163
transform 1 0 33856 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1667941163
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_370
timestamp 1667941163
transform 1 0 35144 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_384
timestamp 1667941163
transform 1 0 36432 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_395
timestamp 1667941163
transform 1 0 37444 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_399
timestamp 1667941163
transform 1 0 37812 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_406
timestamp 1667941163
transform 1 0 38456 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_414
timestamp 1667941163
transform 1 0 39192 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_421
timestamp 1667941163
transform 1 0 39836 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_428
timestamp 1667941163
transform 1 0 40480 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_442
timestamp 1667941163
transform 1 0 41768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_449
timestamp 1667941163
transform 1 0 42412 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_453
timestamp 1667941163
transform 1 0 42780 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_460
timestamp 1667941163
transform 1 0 43424 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_473
timestamp 1667941163
transform 1 0 44620 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_477
timestamp 1667941163
transform 1 0 44988 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_487
timestamp 1667941163
transform 1 0 45908 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_497
timestamp 1667941163
transform 1 0 46828 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_508
timestamp 1667941163
transform 1 0 47840 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_515
timestamp 1667941163
transform 1 0 48484 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_519
timestamp 1667941163
transform 1 0 48852 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_526
timestamp 1667941163
transform 1 0 49496 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_533
timestamp 1667941163
transform 1 0 50140 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_538
timestamp 1667941163
transform 1 0 50600 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_545
timestamp 1667941163
transform 1 0 51244 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_551
timestamp 1667941163
transform 1 0 51796 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_555
timestamp 1667941163
transform 1 0 52164 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_559
timestamp 1667941163
transform 1 0 52532 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_565
timestamp 1667941163
transform 1 0 53084 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_574
timestamp 1667941163
transform 1 0 53912 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_578
timestamp 1667941163
transform 1 0 54280 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_586
timestamp 1667941163
transform 1 0 55016 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_589
timestamp 1667941163
transform 1 0 55292 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_593
timestamp 1667941163
transform 1 0 55660 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_599
timestamp 1667941163
transform 1 0 56212 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_605
timestamp 1667941163
transform 1 0 56764 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_620
timestamp 1667941163
transform 1 0 58144 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_624
timestamp 1667941163
transform 1 0 58512 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1667941163
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1667941163
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1667941163
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_313
timestamp 1667941163
transform 1 0 29900 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_318
timestamp 1667941163
transform 1 0 30360 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_324
timestamp 1667941163
transform 1 0 30912 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_330
timestamp 1667941163
transform 1 0 31464 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1667941163
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_341
timestamp 1667941163
transform 1 0 32476 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_345
timestamp 1667941163
transform 1 0 32844 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_372
timestamp 1667941163
transform 1 0 35328 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_384
timestamp 1667941163
transform 1 0 36432 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_390
timestamp 1667941163
transform 1 0 36984 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_406
timestamp 1667941163
transform 1 0 38456 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_415
timestamp 1667941163
transform 1 0 39284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_429
timestamp 1667941163
transform 1 0 40572 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_433
timestamp 1667941163
transform 1 0 40940 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_442
timestamp 1667941163
transform 1 0 41768 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_449
timestamp 1667941163
transform 1 0 42412 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_455
timestamp 1667941163
transform 1 0 42964 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_462
timestamp 1667941163
transform 1 0 43608 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_466
timestamp 1667941163
transform 1 0 43976 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_488
timestamp 1667941163
transform 1 0 46000 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_492
timestamp 1667941163
transform 1 0 46368 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_500
timestamp 1667941163
transform 1 0 47104 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_505
timestamp 1667941163
transform 1 0 47564 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_515
timestamp 1667941163
transform 1 0 48484 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_530
timestamp 1667941163
transform 1 0 49864 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_536
timestamp 1667941163
transform 1 0 50416 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_544
timestamp 1667941163
transform 1 0 51152 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_555
timestamp 1667941163
transform 1 0 52164 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1667941163
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_561
timestamp 1667941163
transform 1 0 52716 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_567
timestamp 1667941163
transform 1 0 53268 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_576
timestamp 1667941163
transform 1 0 54096 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_584
timestamp 1667941163
transform 1 0 54832 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_592
timestamp 1667941163
transform 1 0 55568 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_603
timestamp 1667941163
transform 1 0 56580 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_613
timestamp 1667941163
transform 1 0 57500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_617
timestamp 1667941163
transform 1 0 57868 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_621
timestamp 1667941163
transform 1 0 58236 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_332
timestamp 1667941163
transform 1 0 31648 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_356
timestamp 1667941163
transform 1 0 33856 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1667941163
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_370
timestamp 1667941163
transform 1 0 35144 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_376
timestamp 1667941163
transform 1 0 35696 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_392
timestamp 1667941163
transform 1 0 37168 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_407
timestamp 1667941163
transform 1 0 38548 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1667941163
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1667941163
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_421
timestamp 1667941163
transform 1 0 39836 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_427
timestamp 1667941163
transform 1 0 40388 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_440
timestamp 1667941163
transform 1 0 41584 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_467
timestamp 1667941163
transform 1 0 44068 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_474
timestamp 1667941163
transform 1 0 44712 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_477
timestamp 1667941163
transform 1 0 44988 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_487
timestamp 1667941163
transform 1 0 45908 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_495
timestamp 1667941163
transform 1 0 46644 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_503
timestamp 1667941163
transform 1 0 47380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_507
timestamp 1667941163
transform 1 0 47748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_512
timestamp 1667941163
transform 1 0 48208 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_520
timestamp 1667941163
transform 1 0 48944 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_526
timestamp 1667941163
transform 1 0 49496 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_533
timestamp 1667941163
transform 1 0 50140 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_538
timestamp 1667941163
transform 1 0 50600 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_544
timestamp 1667941163
transform 1 0 51152 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_550
timestamp 1667941163
transform 1 0 51704 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_558
timestamp 1667941163
transform 1 0 52440 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_562
timestamp 1667941163
transform 1 0 52808 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_570
timestamp 1667941163
transform 1 0 53544 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_582
timestamp 1667941163
transform 1 0 54648 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_589
timestamp 1667941163
transform 1 0 55292 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_599
timestamp 1667941163
transform 1 0 56212 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_603
timestamp 1667941163
transform 1 0 56580 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_611
timestamp 1667941163
transform 1 0 57316 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_623
timestamp 1667941163
transform 1 0 58420 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_302
timestamp 1667941163
transform 1 0 28888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_306
timestamp 1667941163
transform 1 0 29256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_309
timestamp 1667941163
transform 1 0 29532 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_321
timestamp 1667941163
transform 1 0 30636 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_325
timestamp 1667941163
transform 1 0 31004 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_331
timestamp 1667941163
transform 1 0 31556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_360
timestamp 1667941163
transform 1 0 34224 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1667941163
transform 1 0 38180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_412
timestamp 1667941163
transform 1 0 39008 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_428
timestamp 1667941163
transform 1 0 40480 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_51_442
timestamp 1667941163
transform 1 0 41768 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_449
timestamp 1667941163
transform 1 0 42412 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_453
timestamp 1667941163
transform 1 0 42780 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_480
timestamp 1667941163
transform 1 0 45264 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_488
timestamp 1667941163
transform 1 0 46000 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_496
timestamp 1667941163
transform 1 0 46736 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_502
timestamp 1667941163
transform 1 0 47288 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_505
timestamp 1667941163
transform 1 0 47564 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_510
timestamp 1667941163
transform 1 0 48024 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_517
timestamp 1667941163
transform 1 0 48668 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_521
timestamp 1667941163
transform 1 0 49036 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_529
timestamp 1667941163
transform 1 0 49772 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_543
timestamp 1667941163
transform 1 0 51060 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_558
timestamp 1667941163
transform 1 0 52440 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_561
timestamp 1667941163
transform 1 0 52716 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_567
timestamp 1667941163
transform 1 0 53268 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_578
timestamp 1667941163
transform 1 0 54280 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_584
timestamp 1667941163
transform 1 0 54832 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_590
timestamp 1667941163
transform 1 0 55384 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_602
timestamp 1667941163
transform 1 0 56488 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_606
timestamp 1667941163
transform 1 0 56856 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_614
timestamp 1667941163
transform 1 0 57592 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_617
timestamp 1667941163
transform 1 0 57868 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_621
timestamp 1667941163
transform 1 0 58236 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_9
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_335
timestamp 1667941163
transform 1 0 31924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_350
timestamp 1667941163
transform 1 0 33304 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_376
timestamp 1667941163
transform 1 0 35696 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_405
timestamp 1667941163
transform 1 0 38364 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_416
timestamp 1667941163
transform 1 0 39376 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_421
timestamp 1667941163
transform 1 0 39836 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_431
timestamp 1667941163
transform 1 0 40756 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_460
timestamp 1667941163
transform 1 0 43424 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1667941163
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1667941163
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_477
timestamp 1667941163
transform 1 0 44988 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_481
timestamp 1667941163
transform 1 0 45356 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_488
timestamp 1667941163
transform 1 0 46000 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_499
timestamp 1667941163
transform 1 0 47012 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_511
timestamp 1667941163
transform 1 0 48116 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_526
timestamp 1667941163
transform 1 0 49496 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_533
timestamp 1667941163
transform 1 0 50140 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_547
timestamp 1667941163
transform 1 0 51428 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_555
timestamp 1667941163
transform 1 0 52164 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_564
timestamp 1667941163
transform 1 0 52992 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_570
timestamp 1667941163
transform 1 0 53544 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_574
timestamp 1667941163
transform 1 0 53912 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_583
timestamp 1667941163
transform 1 0 54740 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1667941163
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_589
timestamp 1667941163
transform 1 0 55292 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_598
timestamp 1667941163
transform 1 0 56120 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_606
timestamp 1667941163
transform 1 0 56856 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_614
timestamp 1667941163
transform 1 0 57592 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_620
timestamp 1667941163
transform 1 0 58144 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_624
timestamp 1667941163
transform 1 0 58512 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_342
timestamp 1667941163
transform 1 0 32568 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_370
timestamp 1667941163
transform 1 0 35144 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_383
timestamp 1667941163
transform 1 0 36340 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_389
timestamp 1667941163
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_398
timestamp 1667941163
transform 1 0 37720 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_404
timestamp 1667941163
transform 1 0 38272 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_413
timestamp 1667941163
transform 1 0 39100 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_421
timestamp 1667941163
transform 1 0 39836 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_430
timestamp 1667941163
transform 1 0 40664 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_442
timestamp 1667941163
transform 1 0 41768 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_449
timestamp 1667941163
transform 1 0 42412 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_453
timestamp 1667941163
transform 1 0 42780 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_461
timestamp 1667941163
transform 1 0 43516 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_468
timestamp 1667941163
transform 1 0 44160 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_474
timestamp 1667941163
transform 1 0 44712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_481
timestamp 1667941163
transform 1 0 45356 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_494
timestamp 1667941163
transform 1 0 46552 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_501
timestamp 1667941163
transform 1 0 47196 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_505
timestamp 1667941163
transform 1 0 47564 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_512
timestamp 1667941163
transform 1 0 48208 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_525
timestamp 1667941163
transform 1 0 49404 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_533
timestamp 1667941163
transform 1 0 50140 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_542
timestamp 1667941163
transform 1 0 50968 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_552
timestamp 1667941163
transform 1 0 51888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_558
timestamp 1667941163
transform 1 0 52440 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_561
timestamp 1667941163
transform 1 0 52716 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_567
timestamp 1667941163
transform 1 0 53268 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_575
timestamp 1667941163
transform 1 0 54004 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_584
timestamp 1667941163
transform 1 0 54832 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_590
timestamp 1667941163
transform 1 0 55384 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_602
timestamp 1667941163
transform 1 0 56488 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_613
timestamp 1667941163
transform 1 0 57500 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_617
timestamp 1667941163
transform 1 0 57868 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_623
timestamp 1667941163
transform 1 0 58420 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_314
timestamp 1667941163
transform 1 0 29992 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_320
timestamp 1667941163
transform 1 0 30544 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_347
timestamp 1667941163
transform 1 0 33028 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_354
timestamp 1667941163
transform 1 0 33672 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_361
timestamp 1667941163
transform 1 0 34316 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_371
timestamp 1667941163
transform 1 0 35236 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_381
timestamp 1667941163
transform 1 0 36156 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_393
timestamp 1667941163
transform 1 0 37260 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_399
timestamp 1667941163
transform 1 0 37812 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_405
timestamp 1667941163
transform 1 0 38364 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_411
timestamp 1667941163
transform 1 0 38916 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_417
timestamp 1667941163
transform 1 0 39468 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_421
timestamp 1667941163
transform 1 0 39836 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_430
timestamp 1667941163
transform 1 0 40664 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_436
timestamp 1667941163
transform 1 0 41216 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_442
timestamp 1667941163
transform 1 0 41768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_448
timestamp 1667941163
transform 1 0 42320 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_454
timestamp 1667941163
transform 1 0 42872 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_458
timestamp 1667941163
transform 1 0 43240 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_464
timestamp 1667941163
transform 1 0 43792 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_474
timestamp 1667941163
transform 1 0 44712 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_477
timestamp 1667941163
transform 1 0 44988 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_483
timestamp 1667941163
transform 1 0 45540 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_493
timestamp 1667941163
transform 1 0 46460 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_499
timestamp 1667941163
transform 1 0 47012 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_505
timestamp 1667941163
transform 1 0 47564 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_513
timestamp 1667941163
transform 1 0 48300 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_520
timestamp 1667941163
transform 1 0 48944 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_527
timestamp 1667941163
transform 1 0 49588 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1667941163
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_533
timestamp 1667941163
transform 1 0 50140 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_543
timestamp 1667941163
transform 1 0 51060 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_550
timestamp 1667941163
transform 1 0 51704 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_556
timestamp 1667941163
transform 1 0 52256 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_561
timestamp 1667941163
transform 1 0 52716 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_573
timestamp 1667941163
transform 1 0 53820 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_579
timestamp 1667941163
transform 1 0 54372 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_584
timestamp 1667941163
transform 1 0 54832 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_589
timestamp 1667941163
transform 1 0 55292 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_593
timestamp 1667941163
transform 1 0 55660 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_602
timestamp 1667941163
transform 1 0 56488 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_610
timestamp 1667941163
transform 1 0 57224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_618
timestamp 1667941163
transform 1 0 57960 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_624
timestamp 1667941163
transform 1 0 58512 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1667941163
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1667941163
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1667941163
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1667941163
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_319
timestamp 1667941163
transform 1 0 30452 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_326
timestamp 1667941163
transform 1 0 31096 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1667941163
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_342
timestamp 1667941163
transform 1 0 32568 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_366
timestamp 1667941163
transform 1 0 34776 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_378
timestamp 1667941163
transform 1 0 35880 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1667941163
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_397
timestamp 1667941163
transform 1 0 37628 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_409
timestamp 1667941163
transform 1 0 38732 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_421
timestamp 1667941163
transform 1 0 39836 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_432
timestamp 1667941163
transform 1 0 40848 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_443
timestamp 1667941163
transform 1 0 41860 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1667941163
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_449
timestamp 1667941163
transform 1 0 42412 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_458
timestamp 1667941163
transform 1 0 43240 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_462
timestamp 1667941163
transform 1 0 43608 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_484
timestamp 1667941163
transform 1 0 45632 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_490
timestamp 1667941163
transform 1 0 46184 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_496
timestamp 1667941163
transform 1 0 46736 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_502
timestamp 1667941163
transform 1 0 47288 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_505
timestamp 1667941163
transform 1 0 47564 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_513
timestamp 1667941163
transform 1 0 48300 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_521
timestamp 1667941163
transform 1 0 49036 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_529
timestamp 1667941163
transform 1 0 49772 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_535
timestamp 1667941163
transform 1 0 50324 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_544
timestamp 1667941163
transform 1 0 51152 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_556
timestamp 1667941163
transform 1 0 52256 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_561
timestamp 1667941163
transform 1 0 52716 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_571
timestamp 1667941163
transform 1 0 53636 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_585
timestamp 1667941163
transform 1 0 54924 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_591
timestamp 1667941163
transform 1 0 55476 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_600
timestamp 1667941163
transform 1 0 56304 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_611
timestamp 1667941163
transform 1 0 57316 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1667941163
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_617
timestamp 1667941163
transform 1 0 57868 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_621
timestamp 1667941163
transform 1 0 58236 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1667941163
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_314
timestamp 1667941163
transform 1 0 29992 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_318
timestamp 1667941163
transform 1 0 30360 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_322
timestamp 1667941163
transform 1 0 30728 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_349
timestamp 1667941163
transform 1 0 33212 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_356
timestamp 1667941163
transform 1 0 33856 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_371
timestamp 1667941163
transform 1 0 35236 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_381
timestamp 1667941163
transform 1 0 36156 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_388
timestamp 1667941163
transform 1 0 36800 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_399
timestamp 1667941163
transform 1 0 37812 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_405
timestamp 1667941163
transform 1 0 38364 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_414
timestamp 1667941163
transform 1 0 39192 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_56_421
timestamp 1667941163
transform 1 0 39836 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_445
timestamp 1667941163
transform 1 0 42044 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_56_461
timestamp 1667941163
transform 1 0 43516 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_469
timestamp 1667941163
transform 1 0 44252 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_473
timestamp 1667941163
transform 1 0 44620 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_477
timestamp 1667941163
transform 1 0 44988 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_482
timestamp 1667941163
transform 1 0 45448 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_488
timestamp 1667941163
transform 1 0 46000 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_496
timestamp 1667941163
transform 1 0 46736 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_500
timestamp 1667941163
transform 1 0 47104 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_508
timestamp 1667941163
transform 1 0 47840 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_514
timestamp 1667941163
transform 1 0 48392 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_522
timestamp 1667941163
transform 1 0 49128 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_526
timestamp 1667941163
transform 1 0 49496 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_530
timestamp 1667941163
transform 1 0 49864 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_533
timestamp 1667941163
transform 1 0 50140 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_540
timestamp 1667941163
transform 1 0 50784 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_546
timestamp 1667941163
transform 1 0 51336 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_552
timestamp 1667941163
transform 1 0 51888 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_563
timestamp 1667941163
transform 1 0 52900 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_569
timestamp 1667941163
transform 1 0 53452 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_573
timestamp 1667941163
transform 1 0 53820 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1667941163
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1667941163
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_589
timestamp 1667941163
transform 1 0 55292 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_598
timestamp 1667941163
transform 1 0 56120 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_604
timestamp 1667941163
transform 1 0 56672 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_615
timestamp 1667941163
transform 1 0 57684 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_623
timestamp 1667941163
transform 1 0 58420 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_301
timestamp 1667941163
transform 1 0 28796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_307
timestamp 1667941163
transform 1 0 29348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_331
timestamp 1667941163
transform 1 0 31556 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_345
timestamp 1667941163
transform 1 0 32844 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_352
timestamp 1667941163
transform 1 0 33488 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_360
timestamp 1667941163
transform 1 0 34224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_366
timestamp 1667941163
transform 1 0 34776 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_374
timestamp 1667941163
transform 1 0 35512 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_382
timestamp 1667941163
transform 1 0 36248 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1667941163
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_399
timestamp 1667941163
transform 1 0 37812 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_423
timestamp 1667941163
transform 1 0 40020 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_429
timestamp 1667941163
transform 1 0 40572 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_435
timestamp 1667941163
transform 1 0 41124 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_439
timestamp 1667941163
transform 1 0 41492 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_446
timestamp 1667941163
transform 1 0 42136 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_449
timestamp 1667941163
transform 1 0 42412 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_456
timestamp 1667941163
transform 1 0 43056 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_463
timestamp 1667941163
transform 1 0 43700 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_471
timestamp 1667941163
transform 1 0 44436 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_478
timestamp 1667941163
transform 1 0 45080 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_486
timestamp 1667941163
transform 1 0 45816 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_493
timestamp 1667941163
transform 1 0 46460 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_499
timestamp 1667941163
transform 1 0 47012 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1667941163
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_505
timestamp 1667941163
transform 1 0 47564 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_511
timestamp 1667941163
transform 1 0 48116 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_520
timestamp 1667941163
transform 1 0 48944 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_528
timestamp 1667941163
transform 1 0 49680 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_537
timestamp 1667941163
transform 1 0 50508 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_541
timestamp 1667941163
transform 1 0 50876 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_549
timestamp 1667941163
transform 1 0 51612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_558
timestamp 1667941163
transform 1 0 52440 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_561
timestamp 1667941163
transform 1 0 52716 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_571
timestamp 1667941163
transform 1 0 53636 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_581
timestamp 1667941163
transform 1 0 54556 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_587
timestamp 1667941163
transform 1 0 55108 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_593
timestamp 1667941163
transform 1 0 55660 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_599
timestamp 1667941163
transform 1 0 56212 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_607
timestamp 1667941163
transform 1 0 56948 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_614
timestamp 1667941163
transform 1 0 57592 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_617
timestamp 1667941163
transform 1 0 57868 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_621
timestamp 1667941163
transform 1 0 58236 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_285
timestamp 1667941163
transform 1 0 27324 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_297
timestamp 1667941163
transform 1 0 28428 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1667941163
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_331
timestamp 1667941163
transform 1 0 31556 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_341
timestamp 1667941163
transform 1 0 32476 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_356
timestamp 1667941163
transform 1 0 33856 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_387
timestamp 1667941163
transform 1 0 36708 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_400
timestamp 1667941163
transform 1 0 37904 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_404
timestamp 1667941163
transform 1 0 38272 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_411
timestamp 1667941163
transform 1 0 38916 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_418
timestamp 1667941163
transform 1 0 39560 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_421
timestamp 1667941163
transform 1 0 39836 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_425
timestamp 1667941163
transform 1 0 40204 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_449
timestamp 1667941163
transform 1 0 42412 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_459
timestamp 1667941163
transform 1 0 43332 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_474
timestamp 1667941163
transform 1 0 44712 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_477
timestamp 1667941163
transform 1 0 44988 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_481
timestamp 1667941163
transform 1 0 45356 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_491
timestamp 1667941163
transform 1 0 46276 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_504
timestamp 1667941163
transform 1 0 47472 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_510
timestamp 1667941163
transform 1 0 48024 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_521
timestamp 1667941163
transform 1 0 49036 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_528
timestamp 1667941163
transform 1 0 49680 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_533
timestamp 1667941163
transform 1 0 50140 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_539
timestamp 1667941163
transform 1 0 50692 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_548
timestamp 1667941163
transform 1 0 51520 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_555
timestamp 1667941163
transform 1 0 52164 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_563
timestamp 1667941163
transform 1 0 52900 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_570
timestamp 1667941163
transform 1 0 53544 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_576
timestamp 1667941163
transform 1 0 54096 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1667941163
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1667941163
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_589
timestamp 1667941163
transform 1 0 55292 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_593
timestamp 1667941163
transform 1 0 55660 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_601
timestamp 1667941163
transform 1 0 56396 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_607
timestamp 1667941163
transform 1 0 56948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_619
timestamp 1667941163
transform 1 0 58052 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_289
timestamp 1667941163
transform 1 0 27692 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_316
timestamp 1667941163
transform 1 0 30176 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_324
timestamp 1667941163
transform 1 0 30912 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1667941163
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_343
timestamp 1667941163
transform 1 0 32660 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_360
timestamp 1667941163
transform 1 0 34224 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_367
timestamp 1667941163
transform 1 0 34868 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_376
timestamp 1667941163
transform 1 0 35696 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_383
timestamp 1667941163
transform 1 0 36340 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_389
timestamp 1667941163
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_399
timestamp 1667941163
transform 1 0 37812 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_403
timestamp 1667941163
transform 1 0 38180 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_427
timestamp 1667941163
transform 1 0 40388 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_435
timestamp 1667941163
transform 1 0 41124 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_442
timestamp 1667941163
transform 1 0 41768 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_449
timestamp 1667941163
transform 1 0 42412 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_453
timestamp 1667941163
transform 1 0 42780 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_457
timestamp 1667941163
transform 1 0 43148 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_465
timestamp 1667941163
transform 1 0 43884 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_471
timestamp 1667941163
transform 1 0 44436 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_482
timestamp 1667941163
transform 1 0 45448 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_493
timestamp 1667941163
transform 1 0 46460 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_502
timestamp 1667941163
transform 1 0 47288 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_505
timestamp 1667941163
transform 1 0 47564 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_510
timestamp 1667941163
transform 1 0 48024 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_514
timestamp 1667941163
transform 1 0 48392 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_528
timestamp 1667941163
transform 1 0 49680 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_538
timestamp 1667941163
transform 1 0 50600 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_544
timestamp 1667941163
transform 1 0 51152 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_555
timestamp 1667941163
transform 1 0 52164 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1667941163
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_561
timestamp 1667941163
transform 1 0 52716 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_568
timestamp 1667941163
transform 1 0 53360 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_572
timestamp 1667941163
transform 1 0 53728 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_580
timestamp 1667941163
transform 1 0 54464 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_588
timestamp 1667941163
transform 1 0 55200 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_596
timestamp 1667941163
transform 1 0 55936 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_603
timestamp 1667941163
transform 1 0 56580 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_614
timestamp 1667941163
transform 1 0 57592 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_617
timestamp 1667941163
transform 1 0 57868 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_623
timestamp 1667941163
transform 1 0 58420 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_291
timestamp 1667941163
transform 1 0 27876 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_299
timestamp 1667941163
transform 1 0 28612 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_306
timestamp 1667941163
transform 1 0 29256 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_317
timestamp 1667941163
transform 1 0 30268 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_323
timestamp 1667941163
transform 1 0 30820 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_336
timestamp 1667941163
transform 1 0 32016 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_347
timestamp 1667941163
transform 1 0 33028 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_355
timestamp 1667941163
transform 1 0 33764 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_361
timestamp 1667941163
transform 1 0 34316 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_369
timestamp 1667941163
transform 1 0 35052 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_379
timestamp 1667941163
transform 1 0 35972 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_387
timestamp 1667941163
transform 1 0 36708 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_397
timestamp 1667941163
transform 1 0 37628 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_404
timestamp 1667941163
transform 1 0 38272 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_411
timestamp 1667941163
transform 1 0 38916 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_417
timestamp 1667941163
transform 1 0 39468 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_421
timestamp 1667941163
transform 1 0 39836 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_425
timestamp 1667941163
transform 1 0 40204 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_434
timestamp 1667941163
transform 1 0 41032 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_440
timestamp 1667941163
transform 1 0 41584 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_446
timestamp 1667941163
transform 1 0 42136 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_459
timestamp 1667941163
transform 1 0 43332 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_467
timestamp 1667941163
transform 1 0 44068 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_473
timestamp 1667941163
transform 1 0 44620 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_477
timestamp 1667941163
transform 1 0 44988 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_481
timestamp 1667941163
transform 1 0 45356 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_493
timestamp 1667941163
transform 1 0 46460 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_503
timestamp 1667941163
transform 1 0 47380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_509
timestamp 1667941163
transform 1 0 47932 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_515
timestamp 1667941163
transform 1 0 48484 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_524
timestamp 1667941163
transform 1 0 49312 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_530
timestamp 1667941163
transform 1 0 49864 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_533
timestamp 1667941163
transform 1 0 50140 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_548
timestamp 1667941163
transform 1 0 51520 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_556
timestamp 1667941163
transform 1 0 52256 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_560
timestamp 1667941163
transform 1 0 52624 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_563
timestamp 1667941163
transform 1 0 52900 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_569
timestamp 1667941163
transform 1 0 53452 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_574
timestamp 1667941163
transform 1 0 53912 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_580
timestamp 1667941163
transform 1 0 54464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_586
timestamp 1667941163
transform 1 0 55016 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_589
timestamp 1667941163
transform 1 0 55292 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_593
timestamp 1667941163
transform 1 0 55660 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_600
timestamp 1667941163
transform 1 0 56304 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_606
timestamp 1667941163
transform 1 0 56856 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_613
timestamp 1667941163
transform 1 0 57500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_619
timestamp 1667941163
transform 1 0 58052 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_301
timestamp 1667941163
transform 1 0 28796 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_307
timestamp 1667941163
transform 1 0 29348 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_321
timestamp 1667941163
transform 1 0 30636 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_334
timestamp 1667941163
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_346
timestamp 1667941163
transform 1 0 32936 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_363
timestamp 1667941163
transform 1 0 34500 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_378
timestamp 1667941163
transform 1 0 35880 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_399
timestamp 1667941163
transform 1 0 37812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_403
timestamp 1667941163
transform 1 0 38180 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_408
timestamp 1667941163
transform 1 0 38640 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_419
timestamp 1667941163
transform 1 0 39652 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_430
timestamp 1667941163
transform 1 0 40664 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1667941163
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1667941163
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_449
timestamp 1667941163
transform 1 0 42412 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_457
timestamp 1667941163
transform 1 0 43148 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_463
timestamp 1667941163
transform 1 0 43700 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_470
timestamp 1667941163
transform 1 0 44344 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_482
timestamp 1667941163
transform 1 0 45448 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_496
timestamp 1667941163
transform 1 0 46736 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_502
timestamp 1667941163
transform 1 0 47288 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_505
timestamp 1667941163
transform 1 0 47564 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_514
timestamp 1667941163
transform 1 0 48392 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_525
timestamp 1667941163
transform 1 0 49404 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_531
timestamp 1667941163
transform 1 0 49956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_543
timestamp 1667941163
transform 1 0 51060 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_554
timestamp 1667941163
transform 1 0 52072 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_561
timestamp 1667941163
transform 1 0 52716 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_576
timestamp 1667941163
transform 1 0 54096 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_588
timestamp 1667941163
transform 1 0 55200 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_601
timestamp 1667941163
transform 1 0 56396 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_607
timestamp 1667941163
transform 1 0 56948 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_613
timestamp 1667941163
transform 1 0 57500 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_617
timestamp 1667941163
transform 1 0 57868 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_621
timestamp 1667941163
transform 1 0 58236 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1667941163
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_332
timestamp 1667941163
transform 1 0 31648 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_348
timestamp 1667941163
transform 1 0 33120 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_360
timestamp 1667941163
transform 1 0 34224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_373
timestamp 1667941163
transform 1 0 35420 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_379
timestamp 1667941163
transform 1 0 35972 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_387
timestamp 1667941163
transform 1 0 36708 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_393
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_411
timestamp 1667941163
transform 1 0 38916 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_417
timestamp 1667941163
transform 1 0 39468 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_421
timestamp 1667941163
transform 1 0 39836 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_427
timestamp 1667941163
transform 1 0 40388 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_438
timestamp 1667941163
transform 1 0 41400 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_450
timestamp 1667941163
transform 1 0 42504 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_462
timestamp 1667941163
transform 1 0 43608 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_474
timestamp 1667941163
transform 1 0 44712 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_477
timestamp 1667941163
transform 1 0 44988 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_488
timestamp 1667941163
transform 1 0 46000 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_492
timestamp 1667941163
transform 1 0 46368 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_499
timestamp 1667941163
transform 1 0 47012 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_506
timestamp 1667941163
transform 1 0 47656 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_513
timestamp 1667941163
transform 1 0 48300 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_524
timestamp 1667941163
transform 1 0 49312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_530
timestamp 1667941163
transform 1 0 49864 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_533
timestamp 1667941163
transform 1 0 50140 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_543
timestamp 1667941163
transform 1 0 51060 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_547
timestamp 1667941163
transform 1 0 51428 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_550
timestamp 1667941163
transform 1 0 51704 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_558
timestamp 1667941163
transform 1 0 52440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_566
timestamp 1667941163
transform 1 0 53176 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_62_585
timestamp 1667941163
transform 1 0 54924 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_589
timestamp 1667941163
transform 1 0 55292 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_604
timestamp 1667941163
transform 1 0 56672 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_621
timestamp 1667941163
transform 1 0 58236 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1667941163
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1667941163
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1667941163
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1667941163
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_301
timestamp 1667941163
transform 1 0 28796 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_306
timestamp 1667941163
transform 1 0 29256 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_312
timestamp 1667941163
transform 1 0 29808 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1667941163
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_346
timestamp 1667941163
transform 1 0 32936 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_354
timestamp 1667941163
transform 1 0 33672 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_367
timestamp 1667941163
transform 1 0 34868 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_371
timestamp 1667941163
transform 1 0 35236 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_380
timestamp 1667941163
transform 1 0 36064 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_387
timestamp 1667941163
transform 1 0 36708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1667941163
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_399
timestamp 1667941163
transform 1 0 37812 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_407
timestamp 1667941163
transform 1 0 38548 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_414
timestamp 1667941163
transform 1 0 39192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_421
timestamp 1667941163
transform 1 0 39836 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_429
timestamp 1667941163
transform 1 0 40572 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1667941163
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1667941163
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_449
timestamp 1667941163
transform 1 0 42412 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_453
timestamp 1667941163
transform 1 0 42780 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_458
timestamp 1667941163
transform 1 0 43240 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_470
timestamp 1667941163
transform 1 0 44344 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_476
timestamp 1667941163
transform 1 0 44896 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_484
timestamp 1667941163
transform 1 0 45632 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1667941163
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1667941163
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_505
timestamp 1667941163
transform 1 0 47564 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_513
timestamp 1667941163
transform 1 0 48300 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_528
timestamp 1667941163
transform 1 0 49680 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_536
timestamp 1667941163
transform 1 0 50416 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_542
timestamp 1667941163
transform 1 0 50968 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_548
timestamp 1667941163
transform 1 0 51520 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_558
timestamp 1667941163
transform 1 0 52440 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_561
timestamp 1667941163
transform 1 0 52716 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_571
timestamp 1667941163
transform 1 0 53636 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_577
timestamp 1667941163
transform 1 0 54188 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_588
timestamp 1667941163
transform 1 0 55200 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_594
timestamp 1667941163
transform 1 0 55752 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_600
timestamp 1667941163
transform 1 0 56304 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_606
timestamp 1667941163
transform 1 0 56856 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_610
timestamp 1667941163
transform 1 0 57224 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_613
timestamp 1667941163
transform 1 0 57500 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_617
timestamp 1667941163
transform 1 0 57868 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_621
timestamp 1667941163
transform 1 0 58236 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1667941163
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1667941163
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1667941163
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1667941163
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1667941163
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1667941163
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1667941163
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1667941163
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1667941163
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1667941163
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1667941163
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1667941163
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1667941163
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1667941163
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1667941163
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1667941163
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1667941163
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1667941163
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_289
timestamp 1667941163
transform 1 0 27692 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_293
timestamp 1667941163
transform 1 0 28060 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_298
timestamp 1667941163
transform 1 0 28520 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1667941163
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_332
timestamp 1667941163
transform 1 0 31648 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_345
timestamp 1667941163
transform 1 0 32844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_356
timestamp 1667941163
transform 1 0 33856 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1667941163
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_377
timestamp 1667941163
transform 1 0 35788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_389
timestamp 1667941163
transform 1 0 36892 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_395
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_407
timestamp 1667941163
transform 1 0 38548 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_418
timestamp 1667941163
transform 1 0 39560 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_421
timestamp 1667941163
transform 1 0 39836 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_431
timestamp 1667941163
transform 1 0 40756 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_443
timestamp 1667941163
transform 1 0 41860 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_452
timestamp 1667941163
transform 1 0 42688 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_465
timestamp 1667941163
transform 1 0 43884 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_473
timestamp 1667941163
transform 1 0 44620 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_477
timestamp 1667941163
transform 1 0 44988 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_481
timestamp 1667941163
transform 1 0 45356 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_487
timestamp 1667941163
transform 1 0 45908 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_496
timestamp 1667941163
transform 1 0 46736 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_508
timestamp 1667941163
transform 1 0 47840 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_520
timestamp 1667941163
transform 1 0 48944 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_527
timestamp 1667941163
transform 1 0 49588 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1667941163
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_533
timestamp 1667941163
transform 1 0 50140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_537
timestamp 1667941163
transform 1 0 50508 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_551
timestamp 1667941163
transform 1 0 51796 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_557
timestamp 1667941163
transform 1 0 52348 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_563
timestamp 1667941163
transform 1 0 52900 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_567
timestamp 1667941163
transform 1 0 53268 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_572
timestamp 1667941163
transform 1 0 53728 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_584
timestamp 1667941163
transform 1 0 54832 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_589
timestamp 1667941163
transform 1 0 55292 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_602
timestamp 1667941163
transform 1 0 56488 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_614
timestamp 1667941163
transform 1 0 57592 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_619
timestamp 1667941163
transform 1 0 58052 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1667941163
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1667941163
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1667941163
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1667941163
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1667941163
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1667941163
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1667941163
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1667941163
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1667941163
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1667941163
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1667941163
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1667941163
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1667941163
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1667941163
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1667941163
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1667941163
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1667941163
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1667941163
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1667941163
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1667941163
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1667941163
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1667941163
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1667941163
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1667941163
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1667941163
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1667941163
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1667941163
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1667941163
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1667941163
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1667941163
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1667941163
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_293
timestamp 1667941163
transform 1 0 28060 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_301
timestamp 1667941163
transform 1 0 28796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_326
timestamp 1667941163
transform 1 0 31096 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_334
timestamp 1667941163
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_337
timestamp 1667941163
transform 1 0 32108 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_346
timestamp 1667941163
transform 1 0 32936 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_350
timestamp 1667941163
transform 1 0 33304 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_356
timestamp 1667941163
transform 1 0 33856 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_368
timestamp 1667941163
transform 1 0 34960 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_380
timestamp 1667941163
transform 1 0 36064 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_387
timestamp 1667941163
transform 1 0 36708 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1667941163
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_393
timestamp 1667941163
transform 1 0 37260 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_403
timestamp 1667941163
transform 1 0 38180 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_409
timestamp 1667941163
transform 1 0 38732 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_421
timestamp 1667941163
transform 1 0 39836 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_431
timestamp 1667941163
transform 1 0 40756 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1667941163
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1667941163
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_449
timestamp 1667941163
transform 1 0 42412 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_459
timestamp 1667941163
transform 1 0 43332 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_465
timestamp 1667941163
transform 1 0 43884 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_471
timestamp 1667941163
transform 1 0 44436 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_485
timestamp 1667941163
transform 1 0 45724 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_494
timestamp 1667941163
transform 1 0 46552 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_502
timestamp 1667941163
transform 1 0 47288 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_505
timestamp 1667941163
transform 1 0 47564 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_519
timestamp 1667941163
transform 1 0 48852 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_525
timestamp 1667941163
transform 1 0 49404 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_531
timestamp 1667941163
transform 1 0 49956 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_546
timestamp 1667941163
transform 1 0 51336 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_554
timestamp 1667941163
transform 1 0 52072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_558
timestamp 1667941163
transform 1 0 52440 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_561
timestamp 1667941163
transform 1 0 52716 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_576
timestamp 1667941163
transform 1 0 54096 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_582
timestamp 1667941163
transform 1 0 54648 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_588
timestamp 1667941163
transform 1 0 55200 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_601
timestamp 1667941163
transform 1 0 56396 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_612
timestamp 1667941163
transform 1 0 57408 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_617
timestamp 1667941163
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1667941163
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1667941163
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1667941163
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1667941163
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1667941163
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1667941163
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1667941163
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1667941163
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1667941163
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1667941163
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1667941163
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1667941163
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1667941163
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1667941163
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1667941163
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1667941163
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1667941163
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1667941163
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1667941163
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1667941163
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1667941163
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1667941163
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1667941163
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1667941163
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1667941163
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1667941163
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1667941163
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1667941163
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1667941163
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1667941163
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1667941163
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_301
timestamp 1667941163
transform 1 0 28796 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_306
timestamp 1667941163
transform 1 0 29256 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_309
timestamp 1667941163
transform 1 0 29532 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_317
timestamp 1667941163
transform 1 0 30268 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_329
timestamp 1667941163
transform 1 0 31372 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_337
timestamp 1667941163
transform 1 0 32108 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_346
timestamp 1667941163
transform 1 0 32936 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1667941163
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1667941163
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_365
timestamp 1667941163
transform 1 0 34684 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_374
timestamp 1667941163
transform 1 0 35512 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_382
timestamp 1667941163
transform 1 0 36248 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_389
timestamp 1667941163
transform 1 0 36892 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_408
timestamp 1667941163
transform 1 0 38640 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_412
timestamp 1667941163
transform 1 0 39008 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_418
timestamp 1667941163
transform 1 0 39560 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_421
timestamp 1667941163
transform 1 0 39836 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_435
timestamp 1667941163
transform 1 0 41124 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_445
timestamp 1667941163
transform 1 0 42044 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_455
timestamp 1667941163
transform 1 0 42964 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_466
timestamp 1667941163
transform 1 0 43976 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_474
timestamp 1667941163
transform 1 0 44712 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_477
timestamp 1667941163
transform 1 0 44988 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_493
timestamp 1667941163
transform 1 0 46460 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_499
timestamp 1667941163
transform 1 0 47012 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_504
timestamp 1667941163
transform 1 0 47472 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1667941163
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_518
timestamp 1667941163
transform 1 0 48760 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_529
timestamp 1667941163
transform 1 0 49772 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_533
timestamp 1667941163
transform 1 0 50140 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_543
timestamp 1667941163
transform 1 0 51060 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_549
timestamp 1667941163
transform 1 0 51612 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_555
timestamp 1667941163
transform 1 0 52164 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_566
timestamp 1667941163
transform 1 0 53176 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_572
timestamp 1667941163
transform 1 0 53728 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_577
timestamp 1667941163
transform 1 0 54188 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_583
timestamp 1667941163
transform 1 0 54740 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1667941163
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_589
timestamp 1667941163
transform 1 0 55292 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_598
timestamp 1667941163
transform 1 0 56120 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_604
timestamp 1667941163
transform 1 0 56672 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_616
timestamp 1667941163
transform 1 0 57776 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_624
timestamp 1667941163
transform 1 0 58512 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1667941163
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1667941163
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1667941163
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1667941163
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1667941163
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1667941163
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1667941163
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1667941163
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1667941163
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1667941163
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1667941163
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1667941163
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1667941163
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1667941163
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1667941163
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1667941163
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1667941163
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1667941163
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1667941163
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1667941163
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1667941163
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1667941163
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1667941163
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1667941163
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1667941163
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1667941163
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1667941163
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1667941163
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1667941163
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1667941163
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1667941163
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1667941163
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_305
timestamp 1667941163
transform 1 0 29164 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_315
timestamp 1667941163
transform 1 0 30084 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_323
timestamp 1667941163
transform 1 0 30820 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_329
timestamp 1667941163
transform 1 0 31372 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_334
timestamp 1667941163
transform 1 0 31832 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_337
timestamp 1667941163
transform 1 0 32108 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_341
timestamp 1667941163
transform 1 0 32476 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_348
timestamp 1667941163
transform 1 0 33120 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_363
timestamp 1667941163
transform 1 0 34500 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_375
timestamp 1667941163
transform 1 0 35604 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_381
timestamp 1667941163
transform 1 0 36156 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_390
timestamp 1667941163
transform 1 0 36984 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_393
timestamp 1667941163
transform 1 0 37260 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_398
timestamp 1667941163
transform 1 0 37720 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_424
timestamp 1667941163
transform 1 0 40112 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_445
timestamp 1667941163
transform 1 0 42044 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_449
timestamp 1667941163
transform 1 0 42412 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_459
timestamp 1667941163
transform 1 0 43332 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_465
timestamp 1667941163
transform 1 0 43884 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_473
timestamp 1667941163
transform 1 0 44620 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_480
timestamp 1667941163
transform 1 0 45264 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_486
timestamp 1667941163
transform 1 0 45816 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_494
timestamp 1667941163
transform 1 0 46552 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_502
timestamp 1667941163
transform 1 0 47288 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_505
timestamp 1667941163
transform 1 0 47564 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_509
timestamp 1667941163
transform 1 0 47932 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_521
timestamp 1667941163
transform 1 0 49036 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_527
timestamp 1667941163
transform 1 0 49588 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_535
timestamp 1667941163
transform 1 0 50324 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_539
timestamp 1667941163
transform 1 0 50692 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1667941163
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1667941163
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_561
timestamp 1667941163
transform 1 0 52716 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_571
timestamp 1667941163
transform 1 0 53636 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_585
timestamp 1667941163
transform 1 0 54924 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_591
timestamp 1667941163
transform 1 0 55476 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_599
timestamp 1667941163
transform 1 0 56212 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_607
timestamp 1667941163
transform 1 0 56948 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_613
timestamp 1667941163
transform 1 0 57500 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1667941163
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1667941163
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1667941163
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1667941163
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1667941163
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1667941163
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1667941163
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1667941163
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1667941163
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1667941163
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1667941163
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1667941163
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1667941163
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1667941163
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1667941163
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1667941163
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1667941163
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1667941163
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1667941163
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1667941163
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1667941163
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1667941163
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1667941163
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1667941163
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1667941163
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1667941163
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1667941163
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1667941163
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1667941163
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1667941163
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1667941163
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1667941163
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_301
timestamp 1667941163
transform 1 0 28796 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_306
timestamp 1667941163
transform 1 0 29256 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_309
timestamp 1667941163
transform 1 0 29532 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_324
timestamp 1667941163
transform 1 0 30912 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_334
timestamp 1667941163
transform 1 0 31832 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_344
timestamp 1667941163
transform 1 0 32752 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_352
timestamp 1667941163
transform 1 0 33488 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_360
timestamp 1667941163
transform 1 0 34224 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_365
timestamp 1667941163
transform 1 0 34684 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_68_381
timestamp 1667941163
transform 1 0 36156 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_387
timestamp 1667941163
transform 1 0 36708 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_392
timestamp 1667941163
transform 1 0 37168 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_411
timestamp 1667941163
transform 1 0 38916 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_418
timestamp 1667941163
transform 1 0 39560 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_421
timestamp 1667941163
transform 1 0 39836 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_436
timestamp 1667941163
transform 1 0 41216 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_448
timestamp 1667941163
transform 1 0 42320 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_460
timestamp 1667941163
transform 1 0 43424 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_466
timestamp 1667941163
transform 1 0 43976 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_474
timestamp 1667941163
transform 1 0 44712 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_477
timestamp 1667941163
transform 1 0 44988 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_494
timestamp 1667941163
transform 1 0 46552 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_502
timestamp 1667941163
transform 1 0 47288 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_518
timestamp 1667941163
transform 1 0 48760 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_524
timestamp 1667941163
transform 1 0 49312 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_530
timestamp 1667941163
transform 1 0 49864 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_533
timestamp 1667941163
transform 1 0 50140 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_537
timestamp 1667941163
transform 1 0 50508 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_545
timestamp 1667941163
transform 1 0 51244 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_553
timestamp 1667941163
transform 1 0 51980 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_68_561
timestamp 1667941163
transform 1 0 52716 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_571
timestamp 1667941163
transform 1 0 53636 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_583
timestamp 1667941163
transform 1 0 54740 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1667941163
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_589
timestamp 1667941163
transform 1 0 55292 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_599
timestamp 1667941163
transform 1 0 56212 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_620
timestamp 1667941163
transform 1 0 58144 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_624
timestamp 1667941163
transform 1 0 58512 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1667941163
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1667941163
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1667941163
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1667941163
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1667941163
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1667941163
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1667941163
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1667941163
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1667941163
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1667941163
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1667941163
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1667941163
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1667941163
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1667941163
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1667941163
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1667941163
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1667941163
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1667941163
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1667941163
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1667941163
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1667941163
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1667941163
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1667941163
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1667941163
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1667941163
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1667941163
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1667941163
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1667941163
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1667941163
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1667941163
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1667941163
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1667941163
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_305
timestamp 1667941163
transform 1 0 29164 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_313
timestamp 1667941163
transform 1 0 29900 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_318
timestamp 1667941163
transform 1 0 30360 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_330
timestamp 1667941163
transform 1 0 31464 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_69_337
timestamp 1667941163
transform 1 0 32108 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_347
timestamp 1667941163
transform 1 0 33028 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_358
timestamp 1667941163
transform 1 0 34040 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_370
timestamp 1667941163
transform 1 0 35144 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_69_389
timestamp 1667941163
transform 1 0 36892 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_393
timestamp 1667941163
transform 1 0 37260 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_403
timestamp 1667941163
transform 1 0 38180 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_409
timestamp 1667941163
transform 1 0 38732 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_432
timestamp 1667941163
transform 1 0 40848 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_440
timestamp 1667941163
transform 1 0 41584 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_445
timestamp 1667941163
transform 1 0 42044 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_449
timestamp 1667941163
transform 1 0 42412 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_459
timestamp 1667941163
transform 1 0 43332 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_470
timestamp 1667941163
transform 1 0 44344 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_482
timestamp 1667941163
transform 1 0 45448 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_494
timestamp 1667941163
transform 1 0 46552 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_498
timestamp 1667941163
transform 1 0 46920 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_69_505
timestamp 1667941163
transform 1 0 47564 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_509
timestamp 1667941163
transform 1 0 47932 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_513
timestamp 1667941163
transform 1 0 48300 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_521
timestamp 1667941163
transform 1 0 49036 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_532
timestamp 1667941163
transform 1 0 50048 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_540
timestamp 1667941163
transform 1 0 50784 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_547
timestamp 1667941163
transform 1 0 51428 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1667941163
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1667941163
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_561
timestamp 1667941163
transform 1 0 52716 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_568
timestamp 1667941163
transform 1 0 53360 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_576
timestamp 1667941163
transform 1 0 54096 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_582
timestamp 1667941163
transform 1 0 54648 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_590
timestamp 1667941163
transform 1 0 55384 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_596
timestamp 1667941163
transform 1 0 55936 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_602
timestamp 1667941163
transform 1 0 56488 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_610
timestamp 1667941163
transform 1 0 57224 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_69_617
timestamp 1667941163
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1667941163
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1667941163
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1667941163
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1667941163
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1667941163
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1667941163
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1667941163
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1667941163
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1667941163
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1667941163
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1667941163
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1667941163
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1667941163
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1667941163
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1667941163
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1667941163
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1667941163
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1667941163
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1667941163
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1667941163
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1667941163
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1667941163
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1667941163
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1667941163
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1667941163
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1667941163
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1667941163
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1667941163
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1667941163
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1667941163
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_289
timestamp 1667941163
transform 1 0 27692 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_297
timestamp 1667941163
transform 1 0 28428 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_306
timestamp 1667941163
transform 1 0 29256 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_309
timestamp 1667941163
transform 1 0 29532 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_317
timestamp 1667941163
transform 1 0 30268 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_328
timestamp 1667941163
transform 1 0 31280 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_336
timestamp 1667941163
transform 1 0 32016 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_342
timestamp 1667941163
transform 1 0 32568 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_350
timestamp 1667941163
transform 1 0 33304 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_362
timestamp 1667941163
transform 1 0 34408 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_365
timestamp 1667941163
transform 1 0 34684 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_373
timestamp 1667941163
transform 1 0 35420 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_381
timestamp 1667941163
transform 1 0 36156 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_384
timestamp 1667941163
transform 1 0 36432 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_392
timestamp 1667941163
transform 1 0 37168 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_398
timestamp 1667941163
transform 1 0 37720 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_403
timestamp 1667941163
transform 1 0 38180 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_409
timestamp 1667941163
transform 1 0 38732 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_415
timestamp 1667941163
transform 1 0 39284 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1667941163
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_421
timestamp 1667941163
transform 1 0 39836 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_425
timestamp 1667941163
transform 1 0 40204 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_435
timestamp 1667941163
transform 1 0 41124 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_447
timestamp 1667941163
transform 1 0 42228 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_452
timestamp 1667941163
transform 1 0 42688 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_464
timestamp 1667941163
transform 1 0 43792 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_477
timestamp 1667941163
transform 1 0 44988 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_486
timestamp 1667941163
transform 1 0 45816 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_70_505
timestamp 1667941163
transform 1 0 47564 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_70_521
timestamp 1667941163
transform 1 0 49036 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_527
timestamp 1667941163
transform 1 0 49588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_530
timestamp 1667941163
transform 1 0 49864 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_533
timestamp 1667941163
transform 1 0 50140 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_548
timestamp 1667941163
transform 1 0 51520 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_552
timestamp 1667941163
transform 1 0 51888 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_561
timestamp 1667941163
transform 1 0 52716 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_565
timestamp 1667941163
transform 1 0 53084 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_570
timestamp 1667941163
transform 1 0 53544 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_582
timestamp 1667941163
transform 1 0 54648 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_70_589
timestamp 1667941163
transform 1 0 55292 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_604
timestamp 1667941163
transform 1 0 56672 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_608
timestamp 1667941163
transform 1 0 57040 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_622
timestamp 1667941163
transform 1 0 58328 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1667941163
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1667941163
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1667941163
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1667941163
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1667941163
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1667941163
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1667941163
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1667941163
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1667941163
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1667941163
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1667941163
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1667941163
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1667941163
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1667941163
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1667941163
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1667941163
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1667941163
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1667941163
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1667941163
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1667941163
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1667941163
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1667941163
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1667941163
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1667941163
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1667941163
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1667941163
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1667941163
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1667941163
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1667941163
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1667941163
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1667941163
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1667941163
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1667941163
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1667941163
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1667941163
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1667941163
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_337
timestamp 1667941163
transform 1 0 32108 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_346
timestamp 1667941163
transform 1 0 32936 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_357
timestamp 1667941163
transform 1 0 33948 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_369
timestamp 1667941163
transform 1 0 35052 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_379
timestamp 1667941163
transform 1 0 35972 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_387
timestamp 1667941163
transform 1 0 36708 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1667941163
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_393
timestamp 1667941163
transform 1 0 37260 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_399
timestamp 1667941163
transform 1 0 37812 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_411
timestamp 1667941163
transform 1 0 38916 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_417
timestamp 1667941163
transform 1 0 39468 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_425
timestamp 1667941163
transform 1 0 40204 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_431
timestamp 1667941163
transform 1 0 40756 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_439
timestamp 1667941163
transform 1 0 41492 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_446
timestamp 1667941163
transform 1 0 42136 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_449
timestamp 1667941163
transform 1 0 42412 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_459
timestamp 1667941163
transform 1 0 43332 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_470
timestamp 1667941163
transform 1 0 44344 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_482
timestamp 1667941163
transform 1 0 45448 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_488
timestamp 1667941163
transform 1 0 46000 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_502
timestamp 1667941163
transform 1 0 47288 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_505
timestamp 1667941163
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_510
timestamp 1667941163
transform 1 0 48024 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_514
timestamp 1667941163
transform 1 0 48392 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_519
timestamp 1667941163
transform 1 0 48852 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_525
timestamp 1667941163
transform 1 0 49404 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_533
timestamp 1667941163
transform 1 0 50140 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_536
timestamp 1667941163
transform 1 0 50416 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_544
timestamp 1667941163
transform 1 0 51152 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_552
timestamp 1667941163
transform 1 0 51888 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_558
timestamp 1667941163
transform 1 0 52440 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_561
timestamp 1667941163
transform 1 0 52716 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_569
timestamp 1667941163
transform 1 0 53452 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_577
timestamp 1667941163
transform 1 0 54188 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_585
timestamp 1667941163
transform 1 0 54924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_593
timestamp 1667941163
transform 1 0 55660 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_599
timestamp 1667941163
transform 1 0 56212 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_605
timestamp 1667941163
transform 1 0 56764 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_613
timestamp 1667941163
transform 1 0 57500 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1667941163
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1667941163
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1667941163
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1667941163
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1667941163
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1667941163
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1667941163
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1667941163
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1667941163
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1667941163
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1667941163
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1667941163
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1667941163
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1667941163
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1667941163
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1667941163
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1667941163
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1667941163
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1667941163
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1667941163
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1667941163
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1667941163
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1667941163
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1667941163
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1667941163
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1667941163
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1667941163
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1667941163
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1667941163
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1667941163
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1667941163
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_289
timestamp 1667941163
transform 1 0 27692 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_297
timestamp 1667941163
transform 1 0 28428 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_306
timestamp 1667941163
transform 1 0 29256 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_309
timestamp 1667941163
transform 1 0 29532 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_320
timestamp 1667941163
transform 1 0 30544 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_345
timestamp 1667941163
transform 1 0 32844 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_356
timestamp 1667941163
transform 1 0 33856 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_365
timestamp 1667941163
transform 1 0 34684 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_380
timestamp 1667941163
transform 1 0 36064 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_388
timestamp 1667941163
transform 1 0 36800 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_392
timestamp 1667941163
transform 1 0 37168 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_414
timestamp 1667941163
transform 1 0 39192 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_72_421
timestamp 1667941163
transform 1 0 39836 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_432
timestamp 1667941163
transform 1 0 40848 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_442
timestamp 1667941163
transform 1 0 41768 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_72_456
timestamp 1667941163
transform 1 0 43056 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1667941163
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1667941163
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_477
timestamp 1667941163
transform 1 0 44988 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_492
timestamp 1667941163
transform 1 0 46368 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_500
timestamp 1667941163
transform 1 0 47104 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_508
timestamp 1667941163
transform 1 0 47840 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_518
timestamp 1667941163
transform 1 0 48760 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_528
timestamp 1667941163
transform 1 0 49680 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_533
timestamp 1667941163
transform 1 0 50140 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_542
timestamp 1667941163
transform 1 0 50968 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_548
timestamp 1667941163
transform 1 0 51520 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_562
timestamp 1667941163
transform 1 0 52808 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_568
timestamp 1667941163
transform 1 0 53360 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_578
timestamp 1667941163
transform 1 0 54280 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_584
timestamp 1667941163
transform 1 0 54832 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_589
timestamp 1667941163
transform 1 0 55292 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_595
timestamp 1667941163
transform 1 0 55844 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_609
timestamp 1667941163
transform 1 0 57132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_621
timestamp 1667941163
transform 1 0 58236 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1667941163
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1667941163
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1667941163
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1667941163
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1667941163
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1667941163
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1667941163
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1667941163
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1667941163
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1667941163
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1667941163
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1667941163
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1667941163
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1667941163
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1667941163
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1667941163
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1667941163
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1667941163
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1667941163
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1667941163
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1667941163
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1667941163
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1667941163
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1667941163
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1667941163
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1667941163
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1667941163
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1667941163
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1667941163
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1667941163
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1667941163
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1667941163
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_305
timestamp 1667941163
transform 1 0 29164 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_309
timestamp 1667941163
transform 1 0 29532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1667941163
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_329
timestamp 1667941163
transform 1 0 31372 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_334
timestamp 1667941163
transform 1 0 31832 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_337
timestamp 1667941163
transform 1 0 32108 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_345
timestamp 1667941163
transform 1 0 32844 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_357
timestamp 1667941163
transform 1 0 33948 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_360
timestamp 1667941163
transform 1 0 34224 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_368
timestamp 1667941163
transform 1 0 34960 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_374
timestamp 1667941163
transform 1 0 35512 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_377
timestamp 1667941163
transform 1 0 35788 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_387
timestamp 1667941163
transform 1 0 36708 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1667941163
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_393
timestamp 1667941163
transform 1 0 37260 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_399
timestamp 1667941163
transform 1 0 37812 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_405
timestamp 1667941163
transform 1 0 38364 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_416
timestamp 1667941163
transform 1 0 39376 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_422
timestamp 1667941163
transform 1 0 39928 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_426
timestamp 1667941163
transform 1 0 40296 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_434
timestamp 1667941163
transform 1 0 41032 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_446
timestamp 1667941163
transform 1 0 42136 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_449
timestamp 1667941163
transform 1 0 42412 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_455
timestamp 1667941163
transform 1 0 42964 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_467
timestamp 1667941163
transform 1 0 44068 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_473
timestamp 1667941163
transform 1 0 44620 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_484
timestamp 1667941163
transform 1 0 45632 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_496
timestamp 1667941163
transform 1 0 46736 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_502
timestamp 1667941163
transform 1 0 47288 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_505
timestamp 1667941163
transform 1 0 47564 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_515
timestamp 1667941163
transform 1 0 48484 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_529
timestamp 1667941163
transform 1 0 49772 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_535
timestamp 1667941163
transform 1 0 50324 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_546
timestamp 1667941163
transform 1 0 51336 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_552
timestamp 1667941163
transform 1 0 51888 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_558
timestamp 1667941163
transform 1 0 52440 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_561
timestamp 1667941163
transform 1 0 52716 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_567
timestamp 1667941163
transform 1 0 53268 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_575
timestamp 1667941163
transform 1 0 54004 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_584
timestamp 1667941163
transform 1 0 54832 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_590
timestamp 1667941163
transform 1 0 55384 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_596
timestamp 1667941163
transform 1 0 55936 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_602
timestamp 1667941163
transform 1 0 56488 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_614
timestamp 1667941163
transform 1 0 57592 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 1667941163
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1667941163
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1667941163
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1667941163
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1667941163
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1667941163
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1667941163
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1667941163
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1667941163
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1667941163
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1667941163
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1667941163
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1667941163
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1667941163
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1667941163
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1667941163
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1667941163
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1667941163
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1667941163
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1667941163
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1667941163
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1667941163
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1667941163
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1667941163
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1667941163
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1667941163
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1667941163
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1667941163
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1667941163
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1667941163
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1667941163
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1667941163
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1667941163
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1667941163
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1667941163
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_328
timestamp 1667941163
transform 1 0 31280 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_344
timestamp 1667941163
transform 1 0 32752 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_350
timestamp 1667941163
transform 1 0 33304 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_362
timestamp 1667941163
transform 1 0 34408 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_365
timestamp 1667941163
transform 1 0 34684 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_377
timestamp 1667941163
transform 1 0 35788 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_385
timestamp 1667941163
transform 1 0 36524 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_393
timestamp 1667941163
transform 1 0 37260 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_408
timestamp 1667941163
transform 1 0 38640 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_414
timestamp 1667941163
transform 1 0 39192 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_421
timestamp 1667941163
transform 1 0 39836 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_425
timestamp 1667941163
transform 1 0 40204 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_437
timestamp 1667941163
transform 1 0 41308 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_443
timestamp 1667941163
transform 1 0 41860 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_448
timestamp 1667941163
transform 1 0 42320 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_456
timestamp 1667941163
transform 1 0 43056 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_464
timestamp 1667941163
transform 1 0 43792 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_472
timestamp 1667941163
transform 1 0 44528 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_477
timestamp 1667941163
transform 1 0 44988 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_483
timestamp 1667941163
transform 1 0 45540 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_497
timestamp 1667941163
transform 1 0 46828 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_74_507
timestamp 1667941163
transform 1 0 47748 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_513
timestamp 1667941163
transform 1 0 48300 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_518
timestamp 1667941163
transform 1 0 48760 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_530
timestamp 1667941163
transform 1 0 49864 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_533
timestamp 1667941163
transform 1 0 50140 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_537
timestamp 1667941163
transform 1 0 50508 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_543
timestamp 1667941163
transform 1 0 51060 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_74_558
timestamp 1667941163
transform 1 0 52440 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_564
timestamp 1667941163
transform 1 0 52992 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_573
timestamp 1667941163
transform 1 0 53820 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_74_585
timestamp 1667941163
transform 1 0 54924 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_74_589
timestamp 1667941163
transform 1 0 55292 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_602
timestamp 1667941163
transform 1 0 56488 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_606
timestamp 1667941163
transform 1 0 56856 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_620
timestamp 1667941163
transform 1 0 58144 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_624
timestamp 1667941163
transform 1 0 58512 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1667941163
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1667941163
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1667941163
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1667941163
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1667941163
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1667941163
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1667941163
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1667941163
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1667941163
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1667941163
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1667941163
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1667941163
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1667941163
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1667941163
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1667941163
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1667941163
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1667941163
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1667941163
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1667941163
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1667941163
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1667941163
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1667941163
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1667941163
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1667941163
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1667941163
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1667941163
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1667941163
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1667941163
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1667941163
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1667941163
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1667941163
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1667941163
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1667941163
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_317
timestamp 1667941163
transform 1 0 30268 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_327
timestamp 1667941163
transform 1 0 31188 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1667941163
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_337
timestamp 1667941163
transform 1 0 32108 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_343
timestamp 1667941163
transform 1 0 32660 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_351
timestamp 1667941163
transform 1 0 33396 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_362
timestamp 1667941163
transform 1 0 34408 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_75_376
timestamp 1667941163
transform 1 0 35696 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_75_390
timestamp 1667941163
transform 1 0 36984 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_393
timestamp 1667941163
transform 1 0 37260 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_408
timestamp 1667941163
transform 1 0 38640 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_418
timestamp 1667941163
transform 1 0 39560 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_430
timestamp 1667941163
transform 1 0 40664 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_434
timestamp 1667941163
transform 1 0 41032 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_437
timestamp 1667941163
transform 1 0 41308 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_445
timestamp 1667941163
transform 1 0 42044 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_449
timestamp 1667941163
transform 1 0 42412 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_459
timestamp 1667941163
transform 1 0 43332 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_471
timestamp 1667941163
transform 1 0 44436 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_482
timestamp 1667941163
transform 1 0 45448 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_490
timestamp 1667941163
transform 1 0 46184 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_493
timestamp 1667941163
transform 1 0 46460 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_501
timestamp 1667941163
transform 1 0 47196 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_505
timestamp 1667941163
transform 1 0 47564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_509
timestamp 1667941163
transform 1 0 47932 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_514
timestamp 1667941163
transform 1 0 48392 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_522
timestamp 1667941163
transform 1 0 49128 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_75_537
timestamp 1667941163
transform 1 0 50508 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_556
timestamp 1667941163
transform 1 0 52256 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_561
timestamp 1667941163
transform 1 0 52716 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_565
timestamp 1667941163
transform 1 0 53084 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_571
timestamp 1667941163
transform 1 0 53636 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_577
timestamp 1667941163
transform 1 0 54188 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_590
timestamp 1667941163
transform 1 0 55384 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_596
timestamp 1667941163
transform 1 0 55936 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_608
timestamp 1667941163
transform 1 0 57040 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_75_617
timestamp 1667941163
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1667941163
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1667941163
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1667941163
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1667941163
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1667941163
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1667941163
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1667941163
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1667941163
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1667941163
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1667941163
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1667941163
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1667941163
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1667941163
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1667941163
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1667941163
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1667941163
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1667941163
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1667941163
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1667941163
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1667941163
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1667941163
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1667941163
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1667941163
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1667941163
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1667941163
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1667941163
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1667941163
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1667941163
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1667941163
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1667941163
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1667941163
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1667941163
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1667941163
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1667941163
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_321
timestamp 1667941163
transform 1 0 30636 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_329
timestamp 1667941163
transform 1 0 31372 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_344
timestamp 1667941163
transform 1 0 32752 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_354
timestamp 1667941163
transform 1 0 33672 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_360
timestamp 1667941163
transform 1 0 34224 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_365
timestamp 1667941163
transform 1 0 34684 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_369
timestamp 1667941163
transform 1 0 35052 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_373
timestamp 1667941163
transform 1 0 35420 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_376
timestamp 1667941163
transform 1 0 35696 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_386
timestamp 1667941163
transform 1 0 36616 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_396
timestamp 1667941163
transform 1 0 37536 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_412
timestamp 1667941163
transform 1 0 39008 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_418
timestamp 1667941163
transform 1 0 39560 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_421
timestamp 1667941163
transform 1 0 39836 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_434
timestamp 1667941163
transform 1 0 41032 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_442
timestamp 1667941163
transform 1 0 41768 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_454
timestamp 1667941163
transform 1 0 42872 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_462
timestamp 1667941163
transform 1 0 43608 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_468
timestamp 1667941163
transform 1 0 44160 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_474
timestamp 1667941163
transform 1 0 44712 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_477
timestamp 1667941163
transform 1 0 44988 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_486
timestamp 1667941163
transform 1 0 45816 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_490
timestamp 1667941163
transform 1 0 46184 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_493
timestamp 1667941163
transform 1 0 46460 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_505
timestamp 1667941163
transform 1 0 47564 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_517
timestamp 1667941163
transform 1 0 48668 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_528
timestamp 1667941163
transform 1 0 49680 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_533
timestamp 1667941163
transform 1 0 50140 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_543
timestamp 1667941163
transform 1 0 51060 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_553
timestamp 1667941163
transform 1 0 51980 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_559
timestamp 1667941163
transform 1 0 52532 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_565
timestamp 1667941163
transform 1 0 53084 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_576
timestamp 1667941163
transform 1 0 54096 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_582
timestamp 1667941163
transform 1 0 54648 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_76_589
timestamp 1667941163
transform 1 0 55292 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_604
timestamp 1667941163
transform 1 0 56672 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_616
timestamp 1667941163
transform 1 0 57776 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_624
timestamp 1667941163
transform 1 0 58512 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1667941163
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1667941163
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1667941163
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1667941163
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1667941163
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1667941163
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1667941163
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1667941163
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1667941163
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1667941163
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1667941163
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1667941163
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1667941163
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1667941163
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1667941163
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1667941163
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1667941163
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1667941163
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1667941163
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1667941163
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1667941163
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1667941163
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1667941163
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1667941163
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1667941163
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1667941163
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1667941163
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1667941163
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1667941163
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1667941163
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1667941163
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1667941163
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1667941163
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_317
timestamp 1667941163
transform 1 0 30268 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_332
timestamp 1667941163
transform 1 0 31648 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_337
timestamp 1667941163
transform 1 0 32108 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_341
timestamp 1667941163
transform 1 0 32476 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_346
timestamp 1667941163
transform 1 0 32936 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_363
timestamp 1667941163
transform 1 0 34500 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_380
timestamp 1667941163
transform 1 0 36064 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_390
timestamp 1667941163
transform 1 0 36984 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_393
timestamp 1667941163
transform 1 0 37260 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_399
timestamp 1667941163
transform 1 0 37812 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_404
timestamp 1667941163
transform 1 0 38272 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_423
timestamp 1667941163
transform 1 0 40020 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_434
timestamp 1667941163
transform 1 0 41032 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_440
timestamp 1667941163
transform 1 0 41584 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_446
timestamp 1667941163
transform 1 0 42136 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_449
timestamp 1667941163
transform 1 0 42412 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_455
timestamp 1667941163
transform 1 0 42964 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_459
timestamp 1667941163
transform 1 0 43332 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_467
timestamp 1667941163
transform 1 0 44068 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_479
timestamp 1667941163
transform 1 0 45172 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_491
timestamp 1667941163
transform 1 0 46276 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_77_501
timestamp 1667941163
transform 1 0 47196 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_505
timestamp 1667941163
transform 1 0 47564 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_515
timestamp 1667941163
transform 1 0 48484 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_527
timestamp 1667941163
transform 1 0 49588 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_533
timestamp 1667941163
transform 1 0 50140 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_538
timestamp 1667941163
transform 1 0 50600 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_544
timestamp 1667941163
transform 1 0 51152 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_558
timestamp 1667941163
transform 1 0 52440 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_561
timestamp 1667941163
transform 1 0 52716 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_576
timestamp 1667941163
transform 1 0 54096 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_593
timestamp 1667941163
transform 1 0 55660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_605
timestamp 1667941163
transform 1 0 56764 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_613
timestamp 1667941163
transform 1 0 57500 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_617
timestamp 1667941163
transform 1 0 57868 0 -1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1667941163
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1667941163
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1667941163
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1667941163
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1667941163
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1667941163
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1667941163
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1667941163
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1667941163
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1667941163
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1667941163
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1667941163
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1667941163
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1667941163
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1667941163
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1667941163
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1667941163
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1667941163
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1667941163
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1667941163
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1667941163
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1667941163
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1667941163
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1667941163
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1667941163
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1667941163
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1667941163
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1667941163
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1667941163
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1667941163
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1667941163
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1667941163
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1667941163
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1667941163
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_321
timestamp 1667941163
transform 1 0 30636 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_325
timestamp 1667941163
transform 1 0 31004 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_347
timestamp 1667941163
transform 1 0 33028 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_359
timestamp 1667941163
transform 1 0 34132 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1667941163
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_365
timestamp 1667941163
transform 1 0 34684 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_369
timestamp 1667941163
transform 1 0 35052 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_373
timestamp 1667941163
transform 1 0 35420 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_387
timestamp 1667941163
transform 1 0 36708 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_78_414
timestamp 1667941163
transform 1 0 39192 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_421
timestamp 1667941163
transform 1 0 39836 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_425
timestamp 1667941163
transform 1 0 40204 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_431
timestamp 1667941163
transform 1 0 40756 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_435
timestamp 1667941163
transform 1 0 41124 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_442
timestamp 1667941163
transform 1 0 41768 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_454
timestamp 1667941163
transform 1 0 42872 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_465
timestamp 1667941163
transform 1 0 43884 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_471
timestamp 1667941163
transform 1 0 44436 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1667941163
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_477
timestamp 1667941163
transform 1 0 44988 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_492
timestamp 1667941163
transform 1 0 46368 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_502
timestamp 1667941163
transform 1 0 47288 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_508
timestamp 1667941163
transform 1 0 47840 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_519
timestamp 1667941163
transform 1 0 48852 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1667941163
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1667941163
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_533
timestamp 1667941163
transform 1 0 50140 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_542
timestamp 1667941163
transform 1 0 50968 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_78_557
timestamp 1667941163
transform 1 0 52348 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_565
timestamp 1667941163
transform 1 0 53084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_577
timestamp 1667941163
transform 1 0 54188 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_585
timestamp 1667941163
transform 1 0 54924 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1667941163
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1667941163
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1667941163
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1667941163
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1667941163
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1667941163
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1667941163
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1667941163
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1667941163
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1667941163
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1667941163
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1667941163
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1667941163
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1667941163
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1667941163
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1667941163
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1667941163
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1667941163
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1667941163
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1667941163
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1667941163
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1667941163
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1667941163
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1667941163
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1667941163
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1667941163
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1667941163
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1667941163
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1667941163
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1667941163
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1667941163
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1667941163
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1667941163
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1667941163
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1667941163
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1667941163
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_317
timestamp 1667941163
transform 1 0 30268 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_321
timestamp 1667941163
transform 1 0 30636 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1667941163
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1667941163
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_337
timestamp 1667941163
transform 1 0 32108 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_345
timestamp 1667941163
transform 1 0 32844 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_351
timestamp 1667941163
transform 1 0 33396 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_363
timestamp 1667941163
transform 1 0 34500 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_374
timestamp 1667941163
transform 1 0 35512 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_380
timestamp 1667941163
transform 1 0 36064 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_79_390
timestamp 1667941163
transform 1 0 36984 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_393
timestamp 1667941163
transform 1 0 37260 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_397
timestamp 1667941163
transform 1 0 37628 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_408
timestamp 1667941163
transform 1 0 38640 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_414
timestamp 1667941163
transform 1 0 39192 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_422
timestamp 1667941163
transform 1 0 39928 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_434
timestamp 1667941163
transform 1 0 41032 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_446
timestamp 1667941163
transform 1 0 42136 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_449
timestamp 1667941163
transform 1 0 42412 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_453
timestamp 1667941163
transform 1 0 42780 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_461
timestamp 1667941163
transform 1 0 43516 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_469
timestamp 1667941163
transform 1 0 44252 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_79_482
timestamp 1667941163
transform 1 0 45448 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_488
timestamp 1667941163
transform 1 0 46000 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_496
timestamp 1667941163
transform 1 0 46736 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_505
timestamp 1667941163
transform 1 0 47564 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_514
timestamp 1667941163
transform 1 0 48392 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_522
timestamp 1667941163
transform 1 0 49128 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_530
timestamp 1667941163
transform 1 0 49864 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_549
timestamp 1667941163
transform 1 0 51612 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_555
timestamp 1667941163
transform 1 0 52164 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1667941163
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1667941163
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1667941163
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1667941163
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1667941163
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1667941163
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1667941163
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_617
timestamp 1667941163
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1667941163
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1667941163
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1667941163
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1667941163
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1667941163
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1667941163
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1667941163
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1667941163
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1667941163
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1667941163
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1667941163
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1667941163
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1667941163
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1667941163
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1667941163
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1667941163
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1667941163
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1667941163
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1667941163
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1667941163
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1667941163
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1667941163
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1667941163
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1667941163
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1667941163
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1667941163
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1667941163
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1667941163
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1667941163
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1667941163
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1667941163
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1667941163
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1667941163
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1667941163
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_321
timestamp 1667941163
transform 1 0 30636 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_326
timestamp 1667941163
transform 1 0 31096 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_334
timestamp 1667941163
transform 1 0 31832 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_338
timestamp 1667941163
transform 1 0 32200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_347
timestamp 1667941163
transform 1 0 33028 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_355
timestamp 1667941163
transform 1 0 33764 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_361
timestamp 1667941163
transform 1 0 34316 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_80_365
timestamp 1667941163
transform 1 0 34684 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_392
timestamp 1667941163
transform 1 0 37168 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_417
timestamp 1667941163
transform 1 0 39468 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_80_421
timestamp 1667941163
transform 1 0 39836 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_435
timestamp 1667941163
transform 1 0 41124 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_439
timestamp 1667941163
transform 1 0 41492 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_446
timestamp 1667941163
transform 1 0 42136 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_456
timestamp 1667941163
transform 1 0 43056 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_80_470
timestamp 1667941163
transform 1 0 44344 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_80_477
timestamp 1667941163
transform 1 0 44988 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_481
timestamp 1667941163
transform 1 0 45356 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_489
timestamp 1667941163
transform 1 0 46092 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_492
timestamp 1667941163
transform 1 0 46368 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_502
timestamp 1667941163
transform 1 0 47288 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_527
timestamp 1667941163
transform 1 0 49588 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1667941163
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_533
timestamp 1667941163
transform 1 0 50140 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_537
timestamp 1667941163
transform 1 0 50508 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_545
timestamp 1667941163
transform 1 0 51244 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_550
timestamp 1667941163
transform 1 0 51704 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_562
timestamp 1667941163
transform 1 0 52808 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_574
timestamp 1667941163
transform 1 0 53912 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_586
timestamp 1667941163
transform 1 0 55016 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1667941163
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1667941163
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_613
timestamp 1667941163
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1667941163
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1667941163
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1667941163
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1667941163
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1667941163
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1667941163
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1667941163
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1667941163
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1667941163
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1667941163
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1667941163
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1667941163
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1667941163
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1667941163
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1667941163
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1667941163
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1667941163
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1667941163
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1667941163
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1667941163
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1667941163
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1667941163
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1667941163
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1667941163
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1667941163
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1667941163
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1667941163
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1667941163
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1667941163
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1667941163
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1667941163
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1667941163
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1667941163
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_317
timestamp 1667941163
transform 1 0 30268 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_325
timestamp 1667941163
transform 1 0 31004 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_328
timestamp 1667941163
transform 1 0 31280 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_334
timestamp 1667941163
transform 1 0 31832 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_337
timestamp 1667941163
transform 1 0 32108 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_360
timestamp 1667941163
transform 1 0 34224 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1667941163
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1667941163
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_393
timestamp 1667941163
transform 1 0 37260 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_403
timestamp 1667941163
transform 1 0 38180 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_415
timestamp 1667941163
transform 1 0 39284 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_427
timestamp 1667941163
transform 1 0 40388 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_439
timestamp 1667941163
transform 1 0 41492 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_445
timestamp 1667941163
transform 1 0 42044 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_449
timestamp 1667941163
transform 1 0 42412 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_459
timestamp 1667941163
transform 1 0 43332 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_463
timestamp 1667941163
transform 1 0 43700 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_472
timestamp 1667941163
transform 1 0 44528 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_489
timestamp 1667941163
transform 1 0 46092 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_501
timestamp 1667941163
transform 1 0 47196 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_505
timestamp 1667941163
transform 1 0 47564 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_520
timestamp 1667941163
transform 1 0 48944 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_530
timestamp 1667941163
transform 1 0 49864 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_542
timestamp 1667941163
transform 1 0 50968 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_554
timestamp 1667941163
transform 1 0 52072 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1667941163
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1667941163
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1667941163
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1667941163
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1667941163
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1667941163
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1667941163
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1667941163
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1667941163
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1667941163
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1667941163
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1667941163
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1667941163
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1667941163
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1667941163
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1667941163
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1667941163
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1667941163
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1667941163
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1667941163
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1667941163
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1667941163
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1667941163
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1667941163
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1667941163
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1667941163
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1667941163
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1667941163
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1667941163
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1667941163
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1667941163
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1667941163
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1667941163
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1667941163
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1667941163
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1667941163
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1667941163
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1667941163
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1667941163
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1667941163
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1667941163
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1667941163
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_333
timestamp 1667941163
transform 1 0 31740 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_340
timestamp 1667941163
transform 1 0 32384 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_344
timestamp 1667941163
transform 1 0 32752 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_347
timestamp 1667941163
transform 1 0 33028 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_353
timestamp 1667941163
transform 1 0 33580 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_357
timestamp 1667941163
transform 1 0 33948 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_362
timestamp 1667941163
transform 1 0 34408 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_365
timestamp 1667941163
transform 1 0 34684 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_375
timestamp 1667941163
transform 1 0 35604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_381
timestamp 1667941163
transform 1 0 36156 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_385
timestamp 1667941163
transform 1 0 36524 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_390
timestamp 1667941163
transform 1 0 36984 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_398
timestamp 1667941163
transform 1 0 37720 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_403
timestamp 1667941163
transform 1 0 38180 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_411
timestamp 1667941163
transform 1 0 38916 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_417
timestamp 1667941163
transform 1 0 39468 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_421
timestamp 1667941163
transform 1 0 39836 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_427
timestamp 1667941163
transform 1 0 40388 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_435
timestamp 1667941163
transform 1 0 41124 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_441
timestamp 1667941163
transform 1 0 41676 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_456
timestamp 1667941163
transform 1 0 43056 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_462
timestamp 1667941163
transform 1 0 43608 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_468
timestamp 1667941163
transform 1 0 44160 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_474
timestamp 1667941163
transform 1 0 44712 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1667941163
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_486
timestamp 1667941163
transform 1 0 45816 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_497
timestamp 1667941163
transform 1 0 46828 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_509
timestamp 1667941163
transform 1 0 47932 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_521
timestamp 1667941163
transform 1 0 49036 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_529
timestamp 1667941163
transform 1 0 49772 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1667941163
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1667941163
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1667941163
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1667941163
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1667941163
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1667941163
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1667941163
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1667941163
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1667941163
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1667941163
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1667941163
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1667941163
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1667941163
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1667941163
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1667941163
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1667941163
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1667941163
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1667941163
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1667941163
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1667941163
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1667941163
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1667941163
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1667941163
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1667941163
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1667941163
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1667941163
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1667941163
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1667941163
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1667941163
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1667941163
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1667941163
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1667941163
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1667941163
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1667941163
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1667941163
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1667941163
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1667941163
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1667941163
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1667941163
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1667941163
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1667941163
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1667941163
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1667941163
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1667941163
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1667941163
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_337
timestamp 1667941163
transform 1 0 32108 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_346
timestamp 1667941163
transform 1 0 32936 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_357
timestamp 1667941163
transform 1 0 33948 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_83_369
timestamp 1667941163
transform 1 0 35052 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_382
timestamp 1667941163
transform 1 0 36248 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_388
timestamp 1667941163
transform 1 0 36800 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_393
timestamp 1667941163
transform 1 0 37260 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_83_402
timestamp 1667941163
transform 1 0 38088 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_408
timestamp 1667941163
transform 1 0 38640 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_416
timestamp 1667941163
transform 1 0 39376 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_422
timestamp 1667941163
transform 1 0 39928 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_430
timestamp 1667941163
transform 1 0 40664 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_438
timestamp 1667941163
transform 1 0 41400 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_444
timestamp 1667941163
transform 1 0 41952 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_449
timestamp 1667941163
transform 1 0 42412 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_83_458
timestamp 1667941163
transform 1 0 43240 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_466
timestamp 1667941163
transform 1 0 43976 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_83_481
timestamp 1667941163
transform 1 0 45356 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_489
timestamp 1667941163
transform 1 0 46092 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_83_498
timestamp 1667941163
transform 1 0 46920 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1667941163
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1667941163
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1667941163
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1667941163
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1667941163
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1667941163
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1667941163
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1667941163
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1667941163
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1667941163
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1667941163
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1667941163
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_617
timestamp 1667941163
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1667941163
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1667941163
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1667941163
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1667941163
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1667941163
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1667941163
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1667941163
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1667941163
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1667941163
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1667941163
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1667941163
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1667941163
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1667941163
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1667941163
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1667941163
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1667941163
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1667941163
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1667941163
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1667941163
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1667941163
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1667941163
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1667941163
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1667941163
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1667941163
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1667941163
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1667941163
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1667941163
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1667941163
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1667941163
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1667941163
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1667941163
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1667941163
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1667941163
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1667941163
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1667941163
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1667941163
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_84_345
timestamp 1667941163
transform 1 0 32844 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_349
timestamp 1667941163
transform 1 0 33212 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_360
timestamp 1667941163
transform 1 0 34224 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_365
timestamp 1667941163
transform 1 0 34684 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_374
timestamp 1667941163
transform 1 0 35512 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_385
timestamp 1667941163
transform 1 0 36524 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_391
timestamp 1667941163
transform 1 0 37076 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_397
timestamp 1667941163
transform 1 0 37628 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_403
timestamp 1667941163
transform 1 0 38180 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_415
timestamp 1667941163
transform 1 0 39284 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1667941163
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_421
timestamp 1667941163
transform 1 0 39836 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_430
timestamp 1667941163
transform 1 0 40664 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_441
timestamp 1667941163
transform 1 0 41676 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_447
timestamp 1667941163
transform 1 0 42228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_459
timestamp 1667941163
transform 1 0 43332 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_471
timestamp 1667941163
transform 1 0 44436 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1667941163
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1667941163
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1667941163
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1667941163
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1667941163
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1667941163
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1667941163
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1667941163
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1667941163
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1667941163
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1667941163
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1667941163
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1667941163
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1667941163
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1667941163
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1667941163
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1667941163
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1667941163
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1667941163
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1667941163
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1667941163
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1667941163
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1667941163
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1667941163
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1667941163
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1667941163
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1667941163
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1667941163
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1667941163
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1667941163
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1667941163
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1667941163
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1667941163
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1667941163
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1667941163
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1667941163
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1667941163
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1667941163
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1667941163
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1667941163
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1667941163
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1667941163
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1667941163
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1667941163
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1667941163
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1667941163
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1667941163
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1667941163
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1667941163
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1667941163
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1667941163
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1667941163
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1667941163
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_349
timestamp 1667941163
transform 1 0 33212 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_353
timestamp 1667941163
transform 1 0 33580 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_356
timestamp 1667941163
transform 1 0 33856 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_362
timestamp 1667941163
transform 1 0 34408 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_368
timestamp 1667941163
transform 1 0 34960 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_374
timestamp 1667941163
transform 1 0 35512 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_378
timestamp 1667941163
transform 1 0 35880 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_85_386
timestamp 1667941163
transform 1 0 36616 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_85_393
timestamp 1667941163
transform 1 0 37260 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_402
timestamp 1667941163
transform 1 0 38088 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_413
timestamp 1667941163
transform 1 0 39100 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_424
timestamp 1667941163
transform 1 0 40112 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_443
timestamp 1667941163
transform 1 0 41860 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1667941163
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_449
timestamp 1667941163
transform 1 0 42412 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_85_458
timestamp 1667941163
transform 1 0 43240 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_471
timestamp 1667941163
transform 1 0 44436 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_483
timestamp 1667941163
transform 1 0 45540 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_495
timestamp 1667941163
transform 1 0 46644 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1667941163
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1667941163
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1667941163
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1667941163
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1667941163
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1667941163
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1667941163
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1667941163
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1667941163
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1667941163
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1667941163
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1667941163
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1667941163
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_617
timestamp 1667941163
transform 1 0 57868 0 -1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1667941163
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1667941163
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1667941163
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1667941163
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1667941163
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1667941163
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1667941163
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1667941163
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1667941163
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1667941163
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1667941163
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1667941163
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1667941163
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1667941163
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1667941163
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1667941163
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1667941163
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1667941163
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1667941163
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1667941163
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1667941163
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1667941163
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1667941163
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1667941163
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1667941163
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1667941163
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1667941163
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1667941163
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1667941163
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1667941163
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1667941163
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1667941163
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1667941163
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1667941163
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1667941163
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1667941163
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1667941163
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1667941163
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1667941163
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1667941163
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1667941163
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1667941163
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1667941163
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1667941163
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1667941163
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1667941163
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1667941163
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1667941163
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1667941163
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1667941163
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1667941163
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1667941163
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1667941163
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1667941163
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1667941163
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1667941163
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1667941163
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1667941163
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1667941163
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1667941163
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1667941163
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1667941163
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1667941163
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1667941163
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1667941163
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1667941163
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1667941163
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1667941163
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1667941163
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1667941163
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1667941163
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1667941163
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1667941163
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1667941163
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1667941163
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1667941163
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1667941163
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1667941163
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1667941163
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1667941163
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1667941163
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1667941163
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1667941163
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1667941163
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1667941163
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1667941163
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1667941163
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1667941163
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1667941163
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1667941163
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1667941163
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1667941163
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1667941163
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1667941163
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1667941163
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1667941163
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1667941163
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1667941163
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1667941163
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1667941163
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1667941163
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1667941163
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1667941163
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1667941163
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1667941163
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1667941163
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1667941163
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1667941163
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1667941163
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1667941163
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1667941163
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1667941163
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1667941163
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1667941163
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1667941163
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1667941163
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1667941163
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1667941163
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1667941163
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1667941163
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1667941163
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1667941163
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1667941163
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1667941163
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1667941163
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1667941163
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1667941163
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1667941163
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1667941163
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1667941163
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1667941163
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1667941163
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_617
timestamp 1667941163
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1667941163
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1667941163
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1667941163
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1667941163
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1667941163
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1667941163
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1667941163
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1667941163
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1667941163
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1667941163
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1667941163
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1667941163
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1667941163
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1667941163
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1667941163
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1667941163
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1667941163
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1667941163
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1667941163
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1667941163
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1667941163
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1667941163
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1667941163
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1667941163
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1667941163
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1667941163
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1667941163
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1667941163
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1667941163
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1667941163
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1667941163
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1667941163
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1667941163
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1667941163
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1667941163
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1667941163
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1667941163
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1667941163
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1667941163
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1667941163
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1667941163
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1667941163
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1667941163
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1667941163
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1667941163
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1667941163
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1667941163
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1667941163
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1667941163
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1667941163
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1667941163
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1667941163
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1667941163
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1667941163
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1667941163
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1667941163
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1667941163
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1667941163
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1667941163
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1667941163
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1667941163
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1667941163
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1667941163
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1667941163
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1667941163
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1667941163
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1667941163
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1667941163
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1667941163
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1667941163
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1667941163
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1667941163
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1667941163
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1667941163
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1667941163
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1667941163
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1667941163
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1667941163
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1667941163
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1667941163
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1667941163
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1667941163
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1667941163
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1667941163
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1667941163
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1667941163
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1667941163
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1667941163
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1667941163
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1667941163
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1667941163
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1667941163
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1667941163
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1667941163
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1667941163
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1667941163
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1667941163
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1667941163
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1667941163
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1667941163
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1667941163
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1667941163
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1667941163
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1667941163
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1667941163
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1667941163
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1667941163
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1667941163
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1667941163
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1667941163
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1667941163
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1667941163
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1667941163
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1667941163
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1667941163
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1667941163
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1667941163
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1667941163
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1667941163
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1667941163
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1667941163
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1667941163
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1667941163
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1667941163
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1667941163
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1667941163
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1667941163
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1667941163
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1667941163
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1667941163
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1667941163
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1667941163
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1667941163
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1667941163
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1667941163
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1667941163
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1667941163
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1667941163
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1667941163
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1667941163
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1667941163
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1667941163
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1667941163
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1667941163
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1667941163
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1667941163
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1667941163
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1667941163
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1667941163
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1667941163
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1667941163
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1667941163
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1667941163
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1667941163
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1667941163
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1667941163
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1667941163
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1667941163
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1667941163
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1667941163
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1667941163
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1667941163
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1667941163
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1667941163
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1667941163
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1667941163
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1667941163
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1667941163
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1667941163
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1667941163
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1667941163
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1667941163
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1667941163
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1667941163
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1667941163
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1667941163
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1667941163
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1667941163
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1667941163
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1667941163
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1667941163
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1667941163
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1667941163
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1667941163
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1667941163
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1667941163
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1667941163
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1667941163
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1667941163
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1667941163
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1667941163
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1667941163
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1667941163
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1667941163
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1667941163
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1667941163
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1667941163
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1667941163
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_613
timestamp 1667941163
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1667941163
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1667941163
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1667941163
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1667941163
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1667941163
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1667941163
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1667941163
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1667941163
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1667941163
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1667941163
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1667941163
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1667941163
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1667941163
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1667941163
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1667941163
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1667941163
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1667941163
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1667941163
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1667941163
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1667941163
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1667941163
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1667941163
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1667941163
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1667941163
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1667941163
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1667941163
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1667941163
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1667941163
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1667941163
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1667941163
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1667941163
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1667941163
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1667941163
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1667941163
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1667941163
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1667941163
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1667941163
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1667941163
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1667941163
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1667941163
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1667941163
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1667941163
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1667941163
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1667941163
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1667941163
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1667941163
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1667941163
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1667941163
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1667941163
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1667941163
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1667941163
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1667941163
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1667941163
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1667941163
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1667941163
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1667941163
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1667941163
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1667941163
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1667941163
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1667941163
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1667941163
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1667941163
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1667941163
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1667941163
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1667941163
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1667941163
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 1667941163
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1667941163
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1667941163
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1667941163
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1667941163
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1667941163
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1667941163
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1667941163
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1667941163
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1667941163
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1667941163
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1667941163
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1667941163
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1667941163
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1667941163
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1667941163
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1667941163
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1667941163
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1667941163
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1667941163
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1667941163
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1667941163
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1667941163
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1667941163
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1667941163
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1667941163
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1667941163
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1667941163
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1667941163
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1667941163
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1667941163
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1667941163
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1667941163
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1667941163
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1667941163
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1667941163
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1667941163
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1667941163
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1667941163
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1667941163
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1667941163
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1667941163
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1667941163
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1667941163
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1667941163
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1667941163
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1667941163
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1667941163
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1667941163
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1667941163
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1667941163
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1667941163
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1667941163
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1667941163
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1667941163
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1667941163
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1667941163
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1667941163
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1667941163
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1667941163
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1667941163
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1667941163
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1667941163
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1667941163
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1667941163
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1667941163
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1667941163
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1667941163
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1667941163
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1667941163
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1667941163
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1667941163
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1667941163
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1667941163
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1667941163
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1667941163
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1667941163
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1667941163
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1667941163
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1667941163
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1667941163
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1667941163
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1667941163
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1667941163
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1667941163
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1667941163
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1667941163
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1667941163
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1667941163
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1667941163
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1667941163
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1667941163
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1667941163
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1667941163
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1667941163
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1667941163
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1667941163
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1667941163
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1667941163
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1667941163
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1667941163
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1667941163
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1667941163
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1667941163
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1667941163
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1667941163
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1667941163
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1667941163
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1667941163
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1667941163
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1667941163
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1667941163
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1667941163
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1667941163
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1667941163
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1667941163
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1667941163
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1667941163
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1667941163
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1667941163
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1667941163
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1667941163
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1667941163
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1667941163
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1667941163
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1667941163
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1667941163
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1667941163
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1667941163
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1667941163
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1667941163
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1667941163
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1667941163
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_617
timestamp 1667941163
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1667941163
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1667941163
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1667941163
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1667941163
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1667941163
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1667941163
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1667941163
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1667941163
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1667941163
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1667941163
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1667941163
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1667941163
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1667941163
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1667941163
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1667941163
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1667941163
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1667941163
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1667941163
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1667941163
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1667941163
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1667941163
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1667941163
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1667941163
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1667941163
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1667941163
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1667941163
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1667941163
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1667941163
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1667941163
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1667941163
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1667941163
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1667941163
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1667941163
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1667941163
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1667941163
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1667941163
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1667941163
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1667941163
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1667941163
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1667941163
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1667941163
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1667941163
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1667941163
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1667941163
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1667941163
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1667941163
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1667941163
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1667941163
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1667941163
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1667941163
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1667941163
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1667941163
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1667941163
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1667941163
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1667941163
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1667941163
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1667941163
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1667941163
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1667941163
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1667941163
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1667941163
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1667941163
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1667941163
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1667941163
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1667941163
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1667941163
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1667941163
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1667941163
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1667941163
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1667941163
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1667941163
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1667941163
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1667941163
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1667941163
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1667941163
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1667941163
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1667941163
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1667941163
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1667941163
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1667941163
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1667941163
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1667941163
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1667941163
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1667941163
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1667941163
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1667941163
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1667941163
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1667941163
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1667941163
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1667941163
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1667941163
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1667941163
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1667941163
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1667941163
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1667941163
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1667941163
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1667941163
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1667941163
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1667941163
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1667941163
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1667941163
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1667941163
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1667941163
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1667941163
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1667941163
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1667941163
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1667941163
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1667941163
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1667941163
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1667941163
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1667941163
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1667941163
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1667941163
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1667941163
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1667941163
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1667941163
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1667941163
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1667941163
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1667941163
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1667941163
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1667941163
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1667941163
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1667941163
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1667941163
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1667941163
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1667941163
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1667941163
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1667941163
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1667941163
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1667941163
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1667941163
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1667941163
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_617
timestamp 1667941163
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1667941163
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1667941163
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1667941163
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1667941163
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1667941163
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1667941163
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1667941163
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1667941163
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1667941163
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1667941163
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1667941163
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1667941163
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1667941163
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1667941163
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1667941163
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1667941163
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1667941163
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1667941163
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1667941163
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1667941163
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1667941163
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1667941163
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1667941163
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1667941163
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1667941163
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1667941163
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1667941163
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1667941163
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1667941163
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1667941163
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1667941163
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1667941163
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1667941163
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1667941163
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1667941163
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1667941163
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1667941163
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1667941163
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1667941163
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1667941163
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1667941163
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1667941163
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1667941163
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1667941163
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1667941163
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1667941163
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1667941163
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1667941163
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1667941163
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1667941163
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1667941163
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1667941163
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1667941163
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1667941163
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1667941163
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1667941163
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1667941163
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1667941163
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1667941163
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1667941163
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1667941163
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1667941163
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1667941163
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1667941163
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1667941163
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1667941163
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1667941163
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1667941163
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1667941163
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1667941163
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1667941163
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1667941163
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1667941163
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1667941163
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1667941163
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1667941163
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1667941163
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1667941163
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1667941163
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1667941163
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1667941163
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1667941163
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1667941163
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1667941163
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1667941163
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1667941163
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1667941163
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1667941163
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1667941163
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1667941163
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1667941163
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1667941163
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1667941163
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1667941163
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1667941163
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1667941163
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1667941163
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1667941163
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1667941163
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1667941163
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1667941163
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1667941163
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1667941163
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1667941163
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1667941163
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1667941163
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1667941163
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1667941163
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1667941163
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1667941163
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1667941163
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1667941163
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1667941163
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1667941163
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1667941163
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1667941163
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1667941163
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1667941163
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1667941163
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1667941163
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1667941163
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1667941163
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1667941163
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1667941163
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1667941163
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1667941163
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1667941163
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1667941163
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1667941163
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1667941163
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1667941163
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1667941163
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_617
timestamp 1667941163
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1667941163
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1667941163
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1667941163
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1667941163
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1667941163
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1667941163
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1667941163
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1667941163
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1667941163
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1667941163
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1667941163
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1667941163
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1667941163
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1667941163
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1667941163
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1667941163
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1667941163
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1667941163
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1667941163
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1667941163
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1667941163
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1667941163
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1667941163
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1667941163
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1667941163
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1667941163
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1667941163
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1667941163
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1667941163
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1667941163
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1667941163
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1667941163
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1667941163
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1667941163
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1667941163
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1667941163
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1667941163
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1667941163
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1667941163
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1667941163
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1667941163
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1667941163
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1667941163
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1667941163
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1667941163
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1667941163
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1667941163
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1667941163
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1667941163
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1667941163
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1667941163
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1667941163
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1667941163
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1667941163
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1667941163
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1667941163
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1667941163
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1667941163
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1667941163
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1667941163
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1667941163
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1667941163
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1667941163
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1667941163
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1667941163
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1667941163
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_3
timestamp 1667941163
transform 1 0 1380 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_11
timestamp 1667941163
transform 1 0 2116 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_23
timestamp 1667941163
transform 1 0 3220 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_35
timestamp 1667941163
transform 1 0 4324 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_47
timestamp 1667941163
transform 1 0 5428 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1667941163
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1667941163
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1667941163
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1667941163
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1667941163
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1667941163
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1667941163
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1667941163
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1667941163
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1667941163
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1667941163
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1667941163
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1667941163
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1667941163
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1667941163
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1667941163
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1667941163
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1667941163
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1667941163
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1667941163
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1667941163
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1667941163
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1667941163
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1667941163
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1667941163
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1667941163
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1667941163
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1667941163
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1667941163
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1667941163
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1667941163
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1667941163
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1667941163
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1667941163
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1667941163
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1667941163
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1667941163
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1667941163
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1667941163
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1667941163
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1667941163
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1667941163
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1667941163
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1667941163
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1667941163
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1667941163
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1667941163
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1667941163
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1667941163
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1667941163
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1667941163
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1667941163
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1667941163
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1667941163
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1667941163
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1667941163
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1667941163
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1667941163
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1667941163
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1667941163
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1667941163
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_617
timestamp 1667941163
transform 1 0 57868 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_623
timestamp 1667941163
transform 1 0 58420 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_3
timestamp 1667941163
transform 1 0 1380 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_14
timestamp 1667941163
transform 1 0 2392 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_20
timestamp 1667941163
transform 1 0 2944 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1667941163
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1667941163
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1667941163
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1667941163
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1667941163
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1667941163
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1667941163
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1667941163
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1667941163
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1667941163
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1667941163
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1667941163
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1667941163
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1667941163
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1667941163
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1667941163
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1667941163
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1667941163
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1667941163
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1667941163
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1667941163
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1667941163
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1667941163
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1667941163
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1667941163
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1667941163
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1667941163
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1667941163
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1667941163
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1667941163
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1667941163
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1667941163
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1667941163
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1667941163
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1667941163
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1667941163
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1667941163
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1667941163
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1667941163
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1667941163
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1667941163
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1667941163
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1667941163
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1667941163
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1667941163
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1667941163
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1667941163
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1667941163
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1667941163
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1667941163
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1667941163
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1667941163
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1667941163
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1667941163
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1667941163
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1667941163
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1667941163
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1667941163
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1667941163
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1667941163
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1667941163
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1667941163
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_613
timestamp 1667941163
transform 1 0 57500 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_623
timestamp 1667941163
transform 1 0 58420 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_3
timestamp 1667941163
transform 1 0 1380 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_8
timestamp 1667941163
transform 1 0 1840 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_16
timestamp 1667941163
transform 1 0 2576 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_22
timestamp 1667941163
transform 1 0 3128 0 -1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_101_29
timestamp 1667941163
transform 1 0 3772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_41
timestamp 1667941163
transform 1 0 4876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_53
timestamp 1667941163
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1667941163
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1667941163
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_81
timestamp 1667941163
transform 1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_85
timestamp 1667941163
transform 1 0 8924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_97
timestamp 1667941163
transform 1 0 10028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_109
timestamp 1667941163
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1667941163
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1667941163
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_137
timestamp 1667941163
transform 1 0 13708 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_141
timestamp 1667941163
transform 1 0 14076 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_153
timestamp 1667941163
transform 1 0 15180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_165
timestamp 1667941163
transform 1 0 16284 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1667941163
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1667941163
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_193
timestamp 1667941163
transform 1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_197
timestamp 1667941163
transform 1 0 19228 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_209
timestamp 1667941163
transform 1 0 20332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_221
timestamp 1667941163
transform 1 0 21436 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_225
timestamp 1667941163
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1667941163
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_249
timestamp 1667941163
transform 1 0 24012 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_253
timestamp 1667941163
transform 1 0 24380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_265
timestamp 1667941163
transform 1 0 25484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_277
timestamp 1667941163
transform 1 0 26588 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_281
timestamp 1667941163
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_293
timestamp 1667941163
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_305
timestamp 1667941163
transform 1 0 29164 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_309
timestamp 1667941163
transform 1 0 29532 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_321
timestamp 1667941163
transform 1 0 30636 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_333
timestamp 1667941163
transform 1 0 31740 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_337
timestamp 1667941163
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_349
timestamp 1667941163
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_361
timestamp 1667941163
transform 1 0 34316 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_365
timestamp 1667941163
transform 1 0 34684 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_377
timestamp 1667941163
transform 1 0 35788 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_389
timestamp 1667941163
transform 1 0 36892 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_393
timestamp 1667941163
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_405
timestamp 1667941163
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_417
timestamp 1667941163
transform 1 0 39468 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_421
timestamp 1667941163
transform 1 0 39836 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_433
timestamp 1667941163
transform 1 0 40940 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_445
timestamp 1667941163
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1667941163
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1667941163
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_473
timestamp 1667941163
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_477
timestamp 1667941163
transform 1 0 44988 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_489
timestamp 1667941163
transform 1 0 46092 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_501
timestamp 1667941163
transform 1 0 47196 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_505
timestamp 1667941163
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_517
timestamp 1667941163
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_529
timestamp 1667941163
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_533
timestamp 1667941163
transform 1 0 50140 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_545
timestamp 1667941163
transform 1 0 51244 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_557
timestamp 1667941163
transform 1 0 52348 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1667941163
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1667941163
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_585
timestamp 1667941163
transform 1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_589
timestamp 1667941163
transform 1 0 55292 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_601
timestamp 1667941163
transform 1 0 56396 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_613
timestamp 1667941163
transform 1 0 57500 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_617
timestamp 1667941163
transform 1 0 57868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1667941163
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1667941163
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1667941163
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1667941163
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1667941163
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1667941163
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1667941163
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1667941163
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1667941163
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1667941163
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1667941163
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1667941163
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1667941163
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1667941163
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1667941163
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1667941163
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1667941163
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1667941163
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1667941163
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1667941163
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1667941163
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1667941163
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1667941163
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1667941163
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1667941163
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1667941163
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1667941163
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1667941163
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1667941163
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1667941163
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1667941163
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1667941163
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1667941163
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1667941163
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1667941163
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1667941163
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1667941163
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1667941163
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1667941163
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1667941163
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1667941163
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1667941163
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1667941163
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1667941163
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1667941163
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1667941163
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1667941163
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1667941163
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1667941163
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1667941163
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1667941163
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1667941163
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1667941163
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1667941163
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1667941163
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1667941163
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1667941163
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1667941163
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1667941163
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1667941163
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1667941163
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1667941163
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1667941163
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1667941163
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1667941163
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1667941163
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1667941163
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1667941163
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1667941163
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1667941163
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1667941163
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1667941163
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1667941163
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1667941163
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1667941163
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1667941163
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1667941163
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1667941163
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1667941163
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1667941163
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1667941163
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1667941163
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1667941163
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1667941163
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1667941163
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1667941163
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1667941163
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1667941163
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1667941163
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1667941163
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1667941163
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1667941163
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1667941163
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1667941163
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1667941163
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1667941163
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1667941163
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1667941163
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1667941163
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1667941163
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1667941163
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1667941163
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1667941163
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1667941163
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1667941163
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1667941163
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1667941163
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1667941163
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1667941163
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1667941163
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1667941163
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1667941163
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1667941163
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1667941163
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1667941163
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1667941163
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1667941163
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1667941163
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1667941163
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1667941163
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1667941163
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1667941163
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1667941163
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1667941163
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1667941163
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1667941163
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1667941163
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1667941163
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1667941163
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1667941163
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1667941163
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1667941163
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1667941163
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1667941163
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1667941163
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1667941163
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1667941163
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1667941163
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1667941163
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1667941163
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1667941163
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1667941163
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1667941163
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1667941163
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1667941163
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1667941163
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1667941163
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1667941163
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1667941163
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1667941163
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1667941163
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1667941163
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1667941163
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1667941163
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1667941163
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1667941163
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1667941163
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1667941163
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1667941163
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1667941163
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1667941163
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1667941163
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1667941163
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1667941163
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1667941163
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1667941163
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1667941163
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1667941163
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1667941163
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1667941163
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1667941163
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1667941163
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1667941163
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1667941163
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1667941163
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1667941163
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1667941163
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1667941163
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1667941163
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1667941163
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1667941163
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1667941163
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1667941163
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1667941163
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1667941163
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1667941163
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1667941163
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1667941163
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1667941163
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1667941163
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1667941163
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1667941163
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1667941163
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1667941163
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1667941163
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1667941163
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1667941163
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1667941163
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1667941163
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1667941163
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1667941163
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1667941163
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1667941163
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1667941163
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1667941163
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1667941163
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1667941163
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1667941163
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1667941163
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1667941163
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1667941163
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1667941163
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1667941163
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1667941163
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1667941163
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1667941163
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1667941163
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1667941163
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1667941163
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1667941163
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1667941163
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1667941163
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1667941163
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1667941163
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1667941163
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1667941163
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1667941163
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1667941163
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1667941163
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1667941163
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1667941163
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1667941163
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1667941163
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1667941163
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1667941163
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1667941163
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1667941163
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1667941163
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1667941163
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1667941163
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1667941163
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1667941163
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1667941163
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1667941163
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1667941163
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1667941163
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1667941163
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1667941163
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1667941163
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1667941163
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1667941163
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1667941163
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1667941163
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1667941163
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1667941163
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1667941163
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1667941163
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1667941163
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1667941163
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1667941163
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1667941163
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1667941163
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1667941163
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1667941163
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1667941163
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1667941163
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1667941163
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1667941163
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1667941163
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1667941163
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1667941163
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1667941163
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1667941163
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1667941163
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1667941163
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1667941163
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1667941163
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1667941163
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1667941163
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1667941163
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1667941163
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1667941163
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1667941163
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1667941163
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1667941163
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1667941163
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1667941163
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1667941163
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1667941163
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1667941163
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1667941163
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1667941163
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1667941163
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1667941163
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1667941163
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1667941163
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1667941163
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1667941163
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1667941163
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1667941163
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1667941163
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1667941163
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1667941163
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1667941163
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1667941163
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1667941163
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1667941163
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1667941163
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1667941163
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1667941163
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1667941163
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1667941163
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1667941163
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1667941163
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1667941163
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1667941163
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1667941163
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1667941163
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1667941163
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1667941163
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1667941163
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1667941163
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1667941163
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1667941163
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1667941163
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1667941163
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1667941163
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1667941163
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1667941163
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1667941163
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1667941163
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1667941163
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1667941163
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1667941163
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1667941163
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1667941163
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1667941163
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1667941163
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1667941163
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1667941163
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1667941163
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1667941163
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1667941163
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1667941163
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1667941163
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1667941163
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1667941163
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1667941163
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1667941163
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1667941163
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1667941163
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1667941163
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1667941163
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1667941163
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1667941163
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1667941163
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1667941163
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1667941163
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1667941163
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1667941163
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1667941163
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1667941163
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1667941163
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1667941163
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1667941163
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1667941163
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1667941163
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1667941163
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1667941163
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1667941163
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1667941163
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1667941163
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1667941163
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1667941163
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1667941163
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1667941163
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1667941163
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1667941163
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1667941163
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1667941163
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1667941163
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1667941163
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1667941163
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1667941163
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1667941163
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1667941163
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1667941163
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1667941163
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1667941163
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1667941163
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1667941163
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1667941163
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1667941163
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1667941163
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1667941163
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1667941163
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1667941163
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1667941163
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1667941163
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1667941163
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1667941163
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1667941163
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1667941163
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1667941163
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1667941163
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1667941163
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1667941163
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1667941163
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1667941163
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1667941163
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1667941163
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1667941163
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1667941163
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1667941163
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1667941163
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1667941163
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1667941163
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1667941163
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1667941163
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1667941163
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1667941163
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1667941163
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1667941163
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1667941163
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1667941163
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1667941163
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1667941163
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1667941163
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1667941163
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1667941163
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1667941163
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1667941163
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1667941163
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1667941163
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1667941163
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1667941163
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1667941163
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1667941163
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1667941163
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1667941163
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1667941163
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1667941163
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1667941163
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1667941163
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1667941163
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1667941163
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1667941163
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1667941163
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1667941163
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1667941163
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1667941163
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1667941163
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1667941163
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1667941163
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1667941163
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1667941163
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1667941163
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1667941163
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1667941163
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1667941163
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1667941163
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1667941163
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1667941163
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1667941163
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1667941163
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1667941163
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1667941163
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1667941163
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1667941163
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1667941163
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1667941163
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1667941163
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1667941163
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1667941163
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1667941163
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1667941163
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1667941163
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1667941163
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1667941163
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1667941163
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1667941163
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1667941163
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1667941163
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1667941163
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1667941163
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1667941163
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1667941163
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1667941163
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1667941163
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1667941163
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1667941163
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1667941163
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1667941163
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1667941163
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1667941163
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1667941163
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1667941163
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1667941163
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1667941163
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1667941163
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1667941163
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1667941163
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1667941163
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1667941163
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1667941163
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1667941163
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1667941163
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1667941163
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1667941163
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1667941163
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1667941163
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1667941163
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1667941163
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1667941163
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1667941163
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1667941163
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1667941163
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1667941163
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1667941163
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1667941163
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1667941163
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1667941163
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1667941163
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1667941163
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1667941163
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1667941163
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1667941163
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1667941163
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1667941163
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1667941163
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1667941163
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1667941163
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1667941163
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1667941163
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1667941163
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1667941163
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1667941163
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1667941163
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1667941163
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1667941163
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1667941163
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1667941163
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1667941163
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1667941163
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1667941163
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1667941163
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1667941163
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1667941163
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1667941163
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1667941163
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1667941163
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1667941163
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1667941163
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1667941163
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1667941163
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1667941163
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1667941163
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1667941163
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1667941163
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1667941163
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1667941163
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1667941163
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1667941163
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1667941163
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1667941163
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1667941163
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1667941163
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1667941163
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1667941163
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1667941163
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1667941163
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1667941163
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1667941163
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1667941163
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1667941163
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1667941163
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1667941163
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1667941163
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1667941163
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1667941163
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1667941163
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1667941163
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1667941163
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1667941163
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1667941163
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1667941163
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1667941163
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1667941163
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1667941163
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1667941163
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1667941163
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1667941163
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1667941163
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1667941163
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1667941163
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1667941163
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1667941163
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1667941163
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1667941163
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1667941163
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1667941163
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1667941163
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1667941163
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1667941163
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1667941163
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1667941163
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1667941163
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1667941163
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1667941163
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1667941163
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1667941163
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1667941163
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1667941163
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0799_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 46736 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0800_
timestamp 1667941163
transform 1 0 46644 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0801_
timestamp 1667941163
transform -1 0 48116 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0802_
timestamp 1667941163
transform 1 0 48484 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 45172 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0804_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 49956 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0805_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 45908 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0806_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 38456 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a311oi_4  _0807_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 41952 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__or3_1  _0808_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 46460 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0809_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 47564 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0810_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 49312 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform -1 0 48392 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0812_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 47748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0813_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 48760 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0814_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 47012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0815_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 46184 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0816_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 45816 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0817_
timestamp 1667941163
transform 1 0 44252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0818_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 57500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0819_
timestamp 1667941163
transform 1 0 57500 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0820_
timestamp 1667941163
transform -1 0 46552 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0821_
timestamp 1667941163
transform -1 0 46644 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0822_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 38732 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0823_
timestamp 1667941163
transform 1 0 39100 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0824_
timestamp 1667941163
transform -1 0 38364 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0825_
timestamp 1667941163
transform 1 0 36708 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0826_
timestamp 1667941163
transform -1 0 36340 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform -1 0 37720 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0828_
timestamp 1667941163
transform 1 0 36248 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0829_
timestamp 1667941163
transform 1 0 37076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0830_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 40756 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _0831_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 39744 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0832_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0833_
timestamp 1667941163
transform 1 0 38916 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0834_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 42136 0 -1 26112
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0835_
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0836_
timestamp 1667941163
transform -1 0 39284 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0837_
timestamp 1667941163
transform 1 0 40664 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0838_
timestamp 1667941163
transform 1 0 42596 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0839_
timestamp 1667941163
transform -1 0 37444 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0840_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 42596 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0841_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 38180 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0842_
timestamp 1667941163
transform 1 0 38456 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0843_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 38824 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0844_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37444 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0845_
timestamp 1667941163
transform 1 0 36616 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0846_
timestamp 1667941163
transform 1 0 35052 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0847_
timestamp 1667941163
transform -1 0 44712 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0848_
timestamp 1667941163
transform 1 0 45172 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0849_
timestamp 1667941163
transform -1 0 42964 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0850_
timestamp 1667941163
transform 1 0 39100 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0851_
timestamp 1667941163
transform -1 0 41216 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _0852_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0853_
timestamp 1667941163
transform 1 0 38824 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0854_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 42596 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0855_
timestamp 1667941163
transform 1 0 41032 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _0856_
timestamp 1667941163
transform -1 0 38456 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0857_
timestamp 1667941163
transform -1 0 39008 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0858_
timestamp 1667941163
transform 1 0 40020 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0859_
timestamp 1667941163
transform -1 0 45356 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0860_
timestamp 1667941163
transform -1 0 41768 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0861_
timestamp 1667941163
transform 1 0 41492 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0862_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 40664 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0863_
timestamp 1667941163
transform 1 0 39468 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0864_
timestamp 1667941163
transform -1 0 41952 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0865_
timestamp 1667941163
transform 1 0 43884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0866_
timestamp 1667941163
transform 1 0 45908 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0867_
timestamp 1667941163
transform 1 0 40020 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0868_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 38180 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _0869_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 42136 0 -1 27200
box -38 -48 2062 592
use sky130_fd_sc_hd__and3_1  _0870_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 39100 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0871_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 41216 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0872_
timestamp 1667941163
transform 1 0 36708 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0873_
timestamp 1667941163
transform 1 0 39744 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0874_
timestamp 1667941163
transform -1 0 41768 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0875_
timestamp 1667941163
transform 1 0 38456 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0876_
timestamp 1667941163
transform 1 0 40020 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0877_
timestamp 1667941163
transform 1 0 44160 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0878_
timestamp 1667941163
transform -1 0 41768 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0879_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 37996 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0880_
timestamp 1667941163
transform 1 0 35604 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 1667941163
transform 1 0 33580 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0882_
timestamp 1667941163
transform 1 0 35328 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0883_
timestamp 1667941163
transform 1 0 35512 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0884_
timestamp 1667941163
transform 1 0 33672 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0885_
timestamp 1667941163
transform -1 0 40112 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0886_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 39560 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0887_
timestamp 1667941163
transform -1 0 37812 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0888_
timestamp 1667941163
transform -1 0 39192 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0889_
timestamp 1667941163
transform 1 0 35696 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0890_
timestamp 1667941163
transform 1 0 39192 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0891_
timestamp 1667941163
transform -1 0 34776 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0892_
timestamp 1667941163
transform 1 0 36248 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0893_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 37996 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0894_
timestamp 1667941163
transform 1 0 34868 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0895_
timestamp 1667941163
transform -1 0 33304 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0896_
timestamp 1667941163
transform -1 0 38456 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0897_
timestamp 1667941163
transform 1 0 32292 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0898_
timestamp 1667941163
transform -1 0 37812 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0899_
timestamp 1667941163
transform -1 0 37444 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0900_
timestamp 1667941163
transform 1 0 35696 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0901_
timestamp 1667941163
transform -1 0 38916 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0902_
timestamp 1667941163
transform 1 0 31924 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0903_
timestamp 1667941163
transform 1 0 36524 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0904_
timestamp 1667941163
transform 1 0 35788 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0905_
timestamp 1667941163
transform -1 0 35236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0906_
timestamp 1667941163
transform 1 0 40204 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0907_
timestamp 1667941163
transform 1 0 41124 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0908_
timestamp 1667941163
transform 1 0 41492 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0909_
timestamp 1667941163
transform -1 0 41032 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0910_
timestamp 1667941163
transform -1 0 37996 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0911_
timestamp 1667941163
transform 1 0 32292 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0912_
timestamp 1667941163
transform 1 0 40020 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0913_
timestamp 1667941163
transform 1 0 39744 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0914_
timestamp 1667941163
transform -1 0 39100 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0915_
timestamp 1667941163
transform 1 0 29716 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0916_
timestamp 1667941163
transform 1 0 40204 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0917_
timestamp 1667941163
transform 1 0 40020 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0918_
timestamp 1667941163
transform -1 0 29256 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0919_
timestamp 1667941163
transform 1 0 42412 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0920_
timestamp 1667941163
transform 1 0 40756 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0921_
timestamp 1667941163
transform 1 0 28612 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0922_
timestamp 1667941163
transform -1 0 30820 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0923_
timestamp 1667941163
transform -1 0 42044 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0924_
timestamp 1667941163
transform 1 0 38916 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0925_
timestamp 1667941163
transform -1 0 40664 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0926_
timestamp 1667941163
transform 1 0 31280 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0927_
timestamp 1667941163
transform 1 0 40572 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0928_
timestamp 1667941163
transform 1 0 39836 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0929_
timestamp 1667941163
transform 1 0 32292 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0930_
timestamp 1667941163
transform 1 0 41216 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0931_
timestamp 1667941163
transform 1 0 39928 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0932_
timestamp 1667941163
transform 1 0 32292 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0933_
timestamp 1667941163
transform 1 0 36156 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0934_
timestamp 1667941163
transform 1 0 35236 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0935_
timestamp 1667941163
transform 1 0 32568 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0936_
timestamp 1667941163
transform 1 0 33120 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0937_
timestamp 1667941163
transform 1 0 36064 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0938_
timestamp 1667941163
transform 1 0 35328 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 1667941163
transform 1 0 32292 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0940_
timestamp 1667941163
transform -1 0 35052 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0941_
timestamp 1667941163
transform 1 0 36984 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0942_
timestamp 1667941163
transform 1 0 37444 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0943_
timestamp 1667941163
transform 1 0 41584 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0944_
timestamp 1667941163
transform -1 0 41768 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0945_
timestamp 1667941163
transform 1 0 39100 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0946_
timestamp 1667941163
transform 1 0 42504 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0947_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 49312 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0948_
timestamp 1667941163
transform -1 0 36156 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0949_
timestamp 1667941163
transform 1 0 36524 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0950_
timestamp 1667941163
transform 1 0 46736 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0951_
timestamp 1667941163
transform 1 0 49312 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0952_
timestamp 1667941163
transform 1 0 40204 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0953_
timestamp 1667941163
transform 1 0 48116 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0954_
timestamp 1667941163
transform 1 0 48208 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0955_
timestamp 1667941163
transform 1 0 36432 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0956_
timestamp 1667941163
transform -1 0 38916 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0957_
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0958_
timestamp 1667941163
transform -1 0 43424 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0959_
timestamp 1667941163
transform -1 0 41860 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0960_
timestamp 1667941163
transform 1 0 42136 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0961_
timestamp 1667941163
transform 1 0 1564 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0962_
timestamp 1667941163
transform 1 0 1564 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0963_
timestamp 1667941163
transform 1 0 50692 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0964_
timestamp 1667941163
transform -1 0 43148 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1667941163
transform 1 0 42596 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1667941163
transform 1 0 38916 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1667941163
transform 1 0 37444 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1667941163
transform -1 0 41492 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1667941163
transform -1 0 36340 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1667941163
transform 1 0 39284 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1667941163
transform 1 0 32568 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1667941163
transform -1 0 33856 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1667941163
transform 1 0 33028 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1667941163
transform -1 0 32568 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0975_
timestamp 1667941163
transform 1 0 42596 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1667941163
transform 1 0 30084 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1667941163
transform -1 0 29992 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1667941163
transform 1 0 28980 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1667941163
transform -1 0 29992 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1667941163
transform -1 0 31004 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1667941163
transform -1 0 42136 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1667941163
transform 1 0 35420 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1667941163
transform -1 0 30728 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1667941163
transform -1 0 31832 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1667941163
transform -1 0 31096 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0986_
timestamp 1667941163
transform 1 0 43608 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1667941163
transform 1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1667941163
transform -1 0 34316 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1667941163
transform -1 0 35144 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1667941163
transform -1 0 33672 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1667941163
transform 1 0 34132 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1667941163
transform -1 0 44160 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1667941163
transform -1 0 43608 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1667941163
transform 1 0 44344 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1667941163
transform -1 0 43792 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1667941163
transform 1 0 44436 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0997_
timestamp 1667941163
transform -1 0 43056 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1667941163
transform -1 0 43608 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1667941163
transform 1 0 43792 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1000_
timestamp 1667941163
transform 1 0 50600 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1001_
timestamp 1667941163
transform -1 0 35696 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1002_
timestamp 1667941163
transform -1 0 36708 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _1003_
timestamp 1667941163
transform 1 0 35328 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1004_
timestamp 1667941163
transform 1 0 37444 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1005_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34408 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1006_
timestamp 1667941163
transform 1 0 36340 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1007_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34868 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1008_
timestamp 1667941163
transform 1 0 36432 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1009_
timestamp 1667941163
transform -1 0 36248 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1010_
timestamp 1667941163
transform 1 0 36156 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1011_
timestamp 1667941163
transform 1 0 39192 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1012_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 39928 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _1013_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35144 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1014_
timestamp 1667941163
transform 1 0 32476 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1015_
timestamp 1667941163
transform -1 0 36708 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1016_
timestamp 1667941163
transform 1 0 33212 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1017_
timestamp 1667941163
transform -1 0 33120 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1018_
timestamp 1667941163
transform -1 0 33856 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1019_
timestamp 1667941163
transform 1 0 32384 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1020_
timestamp 1667941163
transform -1 0 32844 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1021_
timestamp 1667941163
transform 1 0 32200 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1022_
timestamp 1667941163
transform -1 0 35236 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1023_
timestamp 1667941163
transform -1 0 32568 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1024_
timestamp 1667941163
transform -1 0 38180 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1025_
timestamp 1667941163
transform 1 0 38548 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1026_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 30820 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _1027_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 32936 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1028_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 31832 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  _1029_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32016 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ba_1  _1030_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 31832 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1031_
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1032_
timestamp 1667941163
transform 1 0 30084 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _1033_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 31188 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1034_
timestamp 1667941163
transform 1 0 31464 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1035_
timestamp 1667941163
transform -1 0 33028 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1036_
timestamp 1667941163
transform 1 0 33304 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1037_
timestamp 1667941163
transform -1 0 34500 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _1038_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35236 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__a21oi_1  _1039_
timestamp 1667941163
transform -1 0 36984 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _1040_
timestamp 1667941163
transform 1 0 37536 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _1041_
timestamp 1667941163
transform 1 0 37444 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1042_
timestamp 1667941163
transform 1 0 38732 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1043_
timestamp 1667941163
transform -1 0 38272 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1044_
timestamp 1667941163
transform 1 0 38272 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1045_
timestamp 1667941163
transform -1 0 36984 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _1046_
timestamp 1667941163
transform 1 0 37260 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _1047_
timestamp 1667941163
transform 1 0 37996 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1048_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 38824 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1049_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 40388 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1050_
timestamp 1667941163
transform 1 0 40388 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1051_
timestamp 1667941163
transform 1 0 39560 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1052_
timestamp 1667941163
transform 1 0 40296 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1053_
timestamp 1667941163
transform -1 0 36984 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1054_
timestamp 1667941163
transform 1 0 37444 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1055_
timestamp 1667941163
transform -1 0 33764 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _1056_
timestamp 1667941163
transform 1 0 34592 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _1057_
timestamp 1667941163
transform 1 0 35880 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1058_
timestamp 1667941163
transform 1 0 37444 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1059_
timestamp 1667941163
transform 1 0 40020 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1060_
timestamp 1667941163
transform 1 0 40664 0 -1 48960
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1061_
timestamp 1667941163
transform 1 0 41676 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1062_
timestamp 1667941163
transform -1 0 41676 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _1063_
timestamp 1667941163
transform -1 0 43608 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1064_
timestamp 1667941163
transform 1 0 42872 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1065_
timestamp 1667941163
transform 1 0 39560 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1066_
timestamp 1667941163
transform -1 0 43332 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1067_
timestamp 1667941163
transform -1 0 43332 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1068_
timestamp 1667941163
transform 1 0 43700 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1069_
timestamp 1667941163
transform 1 0 43240 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1070_
timestamp 1667941163
transform 1 0 44068 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1071_
timestamp 1667941163
transform -1 0 46552 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1072_
timestamp 1667941163
transform -1 0 43148 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1073_
timestamp 1667941163
transform 1 0 43240 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1074_
timestamp 1667941163
transform 1 0 40756 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1075_
timestamp 1667941163
transform 1 0 42688 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _1076_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 42504 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1077_
timestamp 1667941163
transform 1 0 41952 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1078_
timestamp 1667941163
transform 1 0 43148 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1079_
timestamp 1667941163
transform 1 0 43608 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1080_
timestamp 1667941163
transform -1 0 41124 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1081_
timestamp 1667941163
transform 1 0 40388 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1082_
timestamp 1667941163
transform 1 0 31004 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _1083_
timestamp 1667941163
transform 1 0 31096 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__o21ai_1  _1084_
timestamp 1667941163
transform -1 0 32384 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1085_
timestamp 1667941163
transform 1 0 32292 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1086_
timestamp 1667941163
transform -1 0 31832 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _1087_
timestamp 1667941163
transform 1 0 32292 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__xor2_1  _1088_
timestamp 1667941163
transform 1 0 32292 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1089_
timestamp 1667941163
transform 1 0 33304 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1090_
timestamp 1667941163
transform 1 0 34040 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1091_
timestamp 1667941163
transform 1 0 34868 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1092_
timestamp 1667941163
transform 1 0 33580 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1093_
timestamp 1667941163
transform 1 0 34868 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1094_
timestamp 1667941163
transform 1 0 35972 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1095_
timestamp 1667941163
transform 1 0 41032 0 1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1096_
timestamp 1667941163
transform 1 0 38548 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1097_
timestamp 1667941163
transform 1 0 39652 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1098_
timestamp 1667941163
transform 1 0 38456 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1099_
timestamp 1667941163
transform 1 0 39468 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1100_
timestamp 1667941163
transform 1 0 42596 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1101_
timestamp 1667941163
transform 1 0 44160 0 -1 47872
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1102_
timestamp 1667941163
transform 1 0 44436 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1103_
timestamp 1667941163
transform -1 0 46552 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1104_
timestamp 1667941163
transform 1 0 48024 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1105_
timestamp 1667941163
transform 1 0 47748 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1106_
timestamp 1667941163
transform 1 0 48760 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1667941163
transform 1 0 44068 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1108_
timestamp 1667941163
transform -1 0 45448 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1109_
timestamp 1667941163
transform 1 0 45172 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1110_
timestamp 1667941163
transform 1 0 45264 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1111_
timestamp 1667941163
transform 1 0 44804 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1112_
timestamp 1667941163
transform 1 0 45816 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1113_
timestamp 1667941163
transform -1 0 44528 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1114_
timestamp 1667941163
transform 1 0 43700 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1115_
timestamp 1667941163
transform 1 0 43792 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1116_
timestamp 1667941163
transform 1 0 44804 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1117_
timestamp 1667941163
transform 1 0 46920 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1667941163
transform 1 0 52256 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1119_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 46460 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1120_
timestamp 1667941163
transform -1 0 47380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1121_
timestamp 1667941163
transform 1 0 32568 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1122_
timestamp 1667941163
transform 1 0 33396 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1123_
timestamp 1667941163
transform -1 0 29256 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _1124_
timestamp 1667941163
transform 1 0 30912 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _1125_
timestamp 1667941163
transform 1 0 31004 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1126_
timestamp 1667941163
transform 1 0 33304 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _1127_
timestamp 1667941163
transform 1 0 34040 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1128_
timestamp 1667941163
transform 1 0 35052 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1129_
timestamp 1667941163
transform 1 0 31464 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1130_
timestamp 1667941163
transform 1 0 32016 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1131_
timestamp 1667941163
transform -1 0 29256 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _1132_
timestamp 1667941163
transform 1 0 29900 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__xor2_1  _1133_
timestamp 1667941163
transform 1 0 30544 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1134_
timestamp 1667941163
transform 1 0 31556 0 1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1135_
timestamp 1667941163
transform 1 0 34868 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1136_
timestamp 1667941163
transform 1 0 35512 0 1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1137_
timestamp 1667941163
transform -1 0 42136 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1138_
timestamp 1667941163
transform 1 0 42596 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1139_
timestamp 1667941163
transform 1 0 40020 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1140_
timestamp 1667941163
transform 1 0 40756 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1141_
timestamp 1667941163
transform 1 0 35604 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1142_
timestamp 1667941163
transform 1 0 40756 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1143_
timestamp 1667941163
transform 1 0 42412 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1144_
timestamp 1667941163
transform 1 0 44896 0 -1 46784
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _1145_
timestamp 1667941163
transform 1 0 41400 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1146_
timestamp 1667941163
transform 1 0 42596 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1147_
timestamp 1667941163
transform 1 0 34592 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1148_
timestamp 1667941163
transform 1 0 34960 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1149_
timestamp 1667941163
transform 1 0 29992 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1150_
timestamp 1667941163
transform 1 0 30728 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1151_
timestamp 1667941163
transform -1 0 29256 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _1152_
timestamp 1667941163
transform 1 0 29164 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__xor2_1  _1153_
timestamp 1667941163
transform 1 0 29624 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1154_
timestamp 1667941163
transform 1 0 30636 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1155_
timestamp 1667941163
transform 1 0 33764 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1156_
timestamp 1667941163
transform 1 0 34868 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1157_
timestamp 1667941163
transform 1 0 43240 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1158_
timestamp 1667941163
transform 1 0 44804 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1159_
timestamp 1667941163
transform -1 0 47012 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1160_
timestamp 1667941163
transform 1 0 46920 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _1161_
timestamp 1667941163
transform -1 0 46736 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1162_
timestamp 1667941163
transform -1 0 47472 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1163_
timestamp 1667941163
transform 1 0 46184 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1164_
timestamp 1667941163
transform -1 0 46552 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1165_
timestamp 1667941163
transform 1 0 46828 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1166_
timestamp 1667941163
transform 1 0 47748 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1167_
timestamp 1667941163
transform 1 0 47748 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1168_
timestamp 1667941163
transform 1 0 48392 0 1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1169_
timestamp 1667941163
transform -1 0 48392 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1170_
timestamp 1667941163
transform 1 0 48852 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1171_
timestamp 1667941163
transform -1 0 37260 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1172_
timestamp 1667941163
transform -1 0 36984 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1173_
timestamp 1667941163
transform 1 0 28888 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1174_
timestamp 1667941163
transform 1 0 30544 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1175_
timestamp 1667941163
transform -1 0 28520 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _1176_
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__xor2_1  _1177_
timestamp 1667941163
transform 1 0 28612 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1178_
timestamp 1667941163
transform 1 0 29900 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1179_
timestamp 1667941163
transform 1 0 32752 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1180_
timestamp 1667941163
transform 1 0 37444 0 -1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1181_
timestamp 1667941163
transform -1 0 42044 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1182_
timestamp 1667941163
transform 1 0 42136 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1183_
timestamp 1667941163
transform 1 0 43424 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1184_
timestamp 1667941163
transform 1 0 45172 0 1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1185_
timestamp 1667941163
transform 1 0 48208 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1186_
timestamp 1667941163
transform 1 0 49036 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1187_
timestamp 1667941163
transform -1 0 49404 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1188_
timestamp 1667941163
transform 1 0 50876 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1189_
timestamp 1667941163
transform 1 0 46828 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1190_
timestamp 1667941163
transform 1 0 49404 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _1191_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 48484 0 -1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_2  _1192_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 49036 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _1193_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 49128 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _1194_
timestamp 1667941163
transform -1 0 49312 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1195_
timestamp 1667941163
transform 1 0 52992 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1196_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 49772 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1197_
timestamp 1667941163
transform 1 0 50324 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1198_
timestamp 1667941163
transform 1 0 50324 0 1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1199_
timestamp 1667941163
transform 1 0 48944 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1200_
timestamp 1667941163
transform -1 0 48024 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _1201_
timestamp 1667941163
transform 1 0 50692 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1202_
timestamp 1667941163
transform -1 0 53268 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1203_
timestamp 1667941163
transform 1 0 49312 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1204_
timestamp 1667941163
transform -1 0 46000 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1205_
timestamp 1667941163
transform -1 0 49496 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1206_
timestamp 1667941163
transform 1 0 51336 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1207_
timestamp 1667941163
transform 1 0 50508 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1208_
timestamp 1667941163
transform -1 0 52164 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1209_
timestamp 1667941163
transform 1 0 52900 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1210_
timestamp 1667941163
transform 1 0 53820 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1211_
timestamp 1667941163
transform 1 0 48484 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1212_
timestamp 1667941163
transform -1 0 49036 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1213_
timestamp 1667941163
transform 1 0 46828 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1214_
timestamp 1667941163
transform -1 0 47564 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1215_
timestamp 1667941163
transform 1 0 43884 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1216_
timestamp 1667941163
transform 1 0 43792 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1217_
timestamp 1667941163
transform 1 0 42596 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1218_
timestamp 1667941163
transform 1 0 45172 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1219_
timestamp 1667941163
transform 1 0 46276 0 -1 47872
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1220_
timestamp 1667941163
transform 1 0 47748 0 -1 46784
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1221_
timestamp 1667941163
transform 1 0 48392 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1222_
timestamp 1667941163
transform 1 0 49404 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1223_
timestamp 1667941163
transform 1 0 46184 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1224_
timestamp 1667941163
transform 1 0 46920 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1225_
timestamp 1667941163
transform -1 0 48484 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1226_
timestamp 1667941163
transform 1 0 47196 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1227_
timestamp 1667941163
transform 1 0 50324 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1228_
timestamp 1667941163
transform 1 0 49220 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1229_
timestamp 1667941163
transform -1 0 48024 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1230_
timestamp 1667941163
transform -1 0 45080 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1231_
timestamp 1667941163
transform 1 0 46644 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1232_
timestamp 1667941163
transform -1 0 46276 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1233_
timestamp 1667941163
transform 1 0 46092 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1234_
timestamp 1667941163
transform 1 0 47196 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1235_
timestamp 1667941163
transform 1 0 47380 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1236_
timestamp 1667941163
transform 1 0 47840 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _1237_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 49496 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1238_
timestamp 1667941163
transform -1 0 49864 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1239_
timestamp 1667941163
transform 1 0 35420 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1240_
timestamp 1667941163
transform -1 0 35880 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1241_
timestamp 1667941163
transform 1 0 38272 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1242_
timestamp 1667941163
transform 1 0 39008 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1243_
timestamp 1667941163
transform 1 0 40020 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1244_
timestamp 1667941163
transform -1 0 38180 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1245_
timestamp 1667941163
transform 1 0 38180 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1246_
timestamp 1667941163
transform -1 0 37812 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _1247_
timestamp 1667941163
transform 1 0 37260 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _1248_
timestamp 1667941163
transform 1 0 37996 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1249_
timestamp 1667941163
transform 1 0 38732 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1250_
timestamp 1667941163
transform 1 0 48208 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1251_
timestamp 1667941163
transform 1 0 34868 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1252_
timestamp 1667941163
transform -1 0 34868 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1253_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37812 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1254_
timestamp 1667941163
transform 1 0 37904 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1255_
timestamp 1667941163
transform 1 0 38916 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1256_
timestamp 1667941163
transform -1 0 37812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1257_
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1258_
timestamp 1667941163
transform -1 0 45908 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1259_
timestamp 1667941163
transform 1 0 45172 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1260_
timestamp 1667941163
transform -1 0 43700 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1261_
timestamp 1667941163
transform -1 0 43056 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1262_
timestamp 1667941163
transform 1 0 42780 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1263_
timestamp 1667941163
transform -1 0 38272 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _1264_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 42780 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1265_
timestamp 1667941163
transform 1 0 45172 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1266_
timestamp 1667941163
transform 1 0 37444 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1267_
timestamp 1667941163
transform -1 0 38916 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1268_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 37628 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1269_
timestamp 1667941163
transform 1 0 37076 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1270_
timestamp 1667941163
transform 1 0 36340 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1271_
timestamp 1667941163
transform -1 0 43240 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1272_
timestamp 1667941163
transform 1 0 43792 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1273_
timestamp 1667941163
transform 1 0 43884 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1274_
timestamp 1667941163
transform 1 0 45172 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1275_
timestamp 1667941163
transform -1 0 45080 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1276_
timestamp 1667941163
transform 1 0 47748 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1277_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 50968 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1278_
timestamp 1667941163
transform 1 0 47012 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1279_
timestamp 1667941163
transform 1 0 48300 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1280_
timestamp 1667941163
transform -1 0 48024 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1281_
timestamp 1667941163
transform -1 0 48024 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1282_
timestamp 1667941163
transform -1 0 51060 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1283_
timestamp 1667941163
transform 1 0 54464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1284_
timestamp 1667941163
transform 1 0 49128 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1285_
timestamp 1667941163
transform -1 0 57224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1286_
timestamp 1667941163
transform 1 0 51428 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1287_
timestamp 1667941163
transform -1 0 52716 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1288_
timestamp 1667941163
transform 1 0 53084 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1289_
timestamp 1667941163
transform 1 0 51612 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1290_
timestamp 1667941163
transform 1 0 51704 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1291_
timestamp 1667941163
transform 1 0 42596 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1292_
timestamp 1667941163
transform 1 0 42136 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1293_
timestamp 1667941163
transform 1 0 39836 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1294_
timestamp 1667941163
transform 1 0 40112 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1295_
timestamp 1667941163
transform -1 0 33304 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1296_
timestamp 1667941163
transform -1 0 33028 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1297_
timestamp 1667941163
transform -1 0 29348 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _1298_
timestamp 1667941163
transform 1 0 29716 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _1299_
timestamp 1667941163
transform 1 0 28612 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1300_
timestamp 1667941163
transform 1 0 32292 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1301_
timestamp 1667941163
transform 1 0 33212 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1302_
timestamp 1667941163
transform 1 0 40388 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1303_
timestamp 1667941163
transform 1 0 45172 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1304_
timestamp 1667941163
transform 1 0 46092 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1305_
timestamp 1667941163
transform 1 0 43424 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1306_
timestamp 1667941163
transform 1 0 43332 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1307_
timestamp 1667941163
transform 1 0 33396 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1308_
timestamp 1667941163
transform 1 0 33488 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _1309_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 34500 0 -1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _1310_
timestamp 1667941163
transform 1 0 29716 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1311_
timestamp 1667941163
transform 1 0 30636 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _1312_
timestamp 1667941163
transform 1 0 29716 0 1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1313_
timestamp 1667941163
transform 1 0 33396 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1314_
timestamp 1667941163
transform 1 0 35052 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1315_
timestamp 1667941163
transform -1 0 35972 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1316_
timestamp 1667941163
transform 1 0 33304 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1317_
timestamp 1667941163
transform 1 0 34868 0 1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1318_
timestamp 1667941163
transform 1 0 44988 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1319_
timestamp 1667941163
transform 1 0 45632 0 1 42432
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1320_
timestamp 1667941163
transform 1 0 51704 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1321_
timestamp 1667941163
transform 1 0 52900 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _1322_
timestamp 1667941163
transform 1 0 52900 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1323_
timestamp 1667941163
transform 1 0 53084 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1324_
timestamp 1667941163
transform 1 0 50232 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1325_
timestamp 1667941163
transform 1 0 50324 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1326_
timestamp 1667941163
transform 1 0 50324 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1327_
timestamp 1667941163
transform 1 0 50416 0 -1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1328_
timestamp 1667941163
transform 1 0 53452 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1329_
timestamp 1667941163
transform 1 0 54464 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _1330_
timestamp 1667941163
transform 1 0 48392 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1331_
timestamp 1667941163
transform 1 0 49128 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1332_
timestamp 1667941163
transform 1 0 49864 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1333_
timestamp 1667941163
transform 1 0 51060 0 -1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1334_
timestamp 1667941163
transform 1 0 53820 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1335_
timestamp 1667941163
transform 1 0 54188 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1336_
timestamp 1667941163
transform 1 0 54004 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1337_
timestamp 1667941163
transform 1 0 49036 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1338_
timestamp 1667941163
transform -1 0 53268 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1339_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 52900 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1340_
timestamp 1667941163
transform 1 0 52256 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1341_
timestamp 1667941163
transform 1 0 51520 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1342_
timestamp 1667941163
transform 1 0 52164 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1343_
timestamp 1667941163
transform 1 0 52900 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1344_
timestamp 1667941163
transform 1 0 49128 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1345_
timestamp 1667941163
transform -1 0 53636 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _1346_
timestamp 1667941163
transform 1 0 53728 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1347_
timestamp 1667941163
transform -1 0 54924 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1348_
timestamp 1667941163
transform -1 0 47288 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1349_
timestamp 1667941163
transform 1 0 48024 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1350_
timestamp 1667941163
transform -1 0 42136 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1351_
timestamp 1667941163
transform 1 0 42320 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1352_
timestamp 1667941163
transform 1 0 35236 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1353_
timestamp 1667941163
transform 1 0 35420 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1354_
timestamp 1667941163
transform -1 0 31832 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1355_
timestamp 1667941163
transform 1 0 32200 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1356_
timestamp 1667941163
transform -1 0 34868 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1357_
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1358_
timestamp 1667941163
transform -1 0 33856 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1359_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33028 0 -1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1360_
timestamp 1667941163
transform 1 0 33304 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1361_
timestamp 1667941163
transform 1 0 33580 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1362_
timestamp 1667941163
transform 1 0 35696 0 -1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1363_
timestamp 1667941163
transform 1 0 43608 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1364_
timestamp 1667941163
transform 1 0 45172 0 1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1365_
timestamp 1667941163
transform 1 0 50692 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1366_
timestamp 1667941163
transform 1 0 51796 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1367_
timestamp 1667941163
transform 1 0 54740 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1368_
timestamp 1667941163
transform 1 0 55476 0 1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__a2bb2o_1  _1369_
timestamp 1667941163
transform -1 0 56304 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1370_
timestamp 1667941163
transform 1 0 55476 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1371_
timestamp 1667941163
transform 1 0 55292 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1372_
timestamp 1667941163
transform -1 0 56580 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1373_
timestamp 1667941163
transform 1 0 55752 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1374_
timestamp 1667941163
transform 1 0 54188 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1375_
timestamp 1667941163
transform -1 0 54556 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1376_
timestamp 1667941163
transform -1 0 37168 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1377_
timestamp 1667941163
transform -1 0 36984 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1378_
timestamp 1667941163
transform 1 0 37444 0 1 38080
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _1379_
timestamp 1667941163
transform 1 0 38088 0 -1 39168
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_1  _1380_
timestamp 1667941163
transform 1 0 33856 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1381_
timestamp 1667941163
transform 1 0 36800 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1382_
timestamp 1667941163
transform 1 0 37444 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1383_
timestamp 1667941163
transform 1 0 37720 0 1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _1384_
timestamp 1667941163
transform 1 0 38824 0 -1 40256
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_1  _1385_
timestamp 1667941163
transform -1 0 42136 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1386_
timestamp 1667941163
transform 1 0 42596 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1387_
timestamp 1667941163
transform 1 0 43700 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1388_
timestamp 1667941163
transform 1 0 46092 0 -1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1389_
timestamp 1667941163
transform 1 0 55016 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1390_
timestamp 1667941163
transform -1 0 51152 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1391_
timestamp 1667941163
transform 1 0 52072 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1392_
timestamp 1667941163
transform 1 0 55936 0 1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _1393_
timestamp 1667941163
transform 1 0 53176 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1394_
timestamp 1667941163
transform 1 0 54096 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1395_
timestamp 1667941163
transform 1 0 55844 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1396_
timestamp 1667941163
transform 1 0 56948 0 1 42432
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1397_
timestamp 1667941163
transform 1 0 56948 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1398_
timestamp 1667941163
transform 1 0 58052 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1399_
timestamp 1667941163
transform 1 0 56948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1400_
timestamp 1667941163
transform 1 0 55752 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1401_
timestamp 1667941163
transform 1 0 52992 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1402_
timestamp 1667941163
transform 1 0 51520 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1403_
timestamp 1667941163
transform 1 0 51980 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _1404_
timestamp 1667941163
transform 1 0 55476 0 1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1405_
timestamp 1667941163
transform 1 0 39100 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1406_
timestamp 1667941163
transform -1 0 39560 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1407_
timestamp 1667941163
transform -1 0 42320 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _1408_
timestamp 1667941163
transform 1 0 40020 0 1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1409_
timestamp 1667941163
transform -1 0 42044 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1410_
timestamp 1667941163
transform 1 0 42596 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1411_
timestamp 1667941163
transform -1 0 36892 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _1412_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 36708 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1413_
timestamp 1667941163
transform 1 0 36248 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1414_
timestamp 1667941163
transform -1 0 36064 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1415_
timestamp 1667941163
transform -1 0 36892 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1416_
timestamp 1667941163
transform 1 0 43700 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1417_
timestamp 1667941163
transform 1 0 45172 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1418_
timestamp 1667941163
transform 1 0 46368 0 1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _1419_
timestamp 1667941163
transform 1 0 53728 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1420_
timestamp 1667941163
transform 1 0 53912 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1421_
timestamp 1667941163
transform 1 0 54740 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1422_
timestamp 1667941163
transform 1 0 56580 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1423_
timestamp 1667941163
transform 1 0 57132 0 1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__a2bb2o_1  _1424_
timestamp 1667941163
transform -1 0 56488 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1425_
timestamp 1667941163
transform -1 0 57316 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1426_
timestamp 1667941163
transform 1 0 57040 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _1427_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 57040 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1428_
timestamp 1667941163
transform -1 0 58420 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1429_
timestamp 1667941163
transform -1 0 56488 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1430_
timestamp 1667941163
transform -1 0 57500 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1431_
timestamp 1667941163
transform -1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1432_
timestamp 1667941163
transform 1 0 48300 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1433_
timestamp 1667941163
transform 1 0 39468 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1434_
timestamp 1667941163
transform 1 0 40388 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1435_
timestamp 1667941163
transform 1 0 40848 0 -1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1436_
timestamp 1667941163
transform -1 0 42688 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1437_
timestamp 1667941163
transform 1 0 42688 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1438_
timestamp 1667941163
transform 1 0 44068 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1439_
timestamp 1667941163
transform 1 0 45356 0 1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1440_
timestamp 1667941163
transform 1 0 55568 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1441_
timestamp 1667941163
transform 1 0 53268 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1442_
timestamp 1667941163
transform 1 0 54004 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1443_
timestamp 1667941163
transform 1 0 56304 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1444_
timestamp 1667941163
transform 1 0 56948 0 1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1445_
timestamp 1667941163
transform 1 0 56948 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1446_
timestamp 1667941163
transform -1 0 57960 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1447_
timestamp 1667941163
transform -1 0 58420 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1448_
timestamp 1667941163
transform -1 0 39192 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1449_
timestamp 1667941163
transform -1 0 38180 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1450_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 40756 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1451_
timestamp 1667941163
transform 1 0 43332 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1452_
timestamp 1667941163
transform 1 0 42228 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1453_
timestamp 1667941163
transform 1 0 44988 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1454_
timestamp 1667941163
transform 1 0 42596 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1455_
timestamp 1667941163
transform 1 0 43976 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1456_
timestamp 1667941163
transform 1 0 45264 0 1 38080
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1457_
timestamp 1667941163
transform 1 0 51612 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1458_
timestamp 1667941163
transform -1 0 53636 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1459_
timestamp 1667941163
transform 1 0 52532 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1460_
timestamp 1667941163
transform 1 0 55844 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1461_
timestamp 1667941163
transform 1 0 53820 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1462_
timestamp 1667941163
transform 1 0 54188 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1463_
timestamp 1667941163
transform 1 0 55476 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1464_
timestamp 1667941163
transform 1 0 56764 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1465_
timestamp 1667941163
transform 1 0 54004 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1466_
timestamp 1667941163
transform -1 0 54280 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1467_
timestamp 1667941163
transform 1 0 55752 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1468_
timestamp 1667941163
transform -1 0 47288 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1469_
timestamp 1667941163
transform 1 0 48116 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1470_
timestamp 1667941163
transform 1 0 41492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1471_
timestamp 1667941163
transform 1 0 42596 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1472_
timestamp 1667941163
transform 1 0 43240 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1473_
timestamp 1667941163
transform 1 0 44528 0 -1 38080
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1474_
timestamp 1667941163
transform 1 0 50692 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1475_
timestamp 1667941163
transform 1 0 52900 0 -1 38080
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _1476_
timestamp 1667941163
transform -1 0 53912 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1477_
timestamp 1667941163
transform 1 0 54464 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1478_
timestamp 1667941163
transform 1 0 55752 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1479_
timestamp 1667941163
transform -1 0 58236 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1480_
timestamp 1667941163
transform 1 0 56672 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1481_
timestamp 1667941163
transform -1 0 54832 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1482_
timestamp 1667941163
transform -1 0 56120 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1483_
timestamp 1667941163
transform 1 0 56948 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1484_
timestamp 1667941163
transform 1 0 57316 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1485_
timestamp 1667941163
transform 1 0 56948 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1486_
timestamp 1667941163
transform -1 0 58420 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1487_
timestamp 1667941163
transform 1 0 57224 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1488_
timestamp 1667941163
transform 1 0 48760 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1489_
timestamp 1667941163
transform -1 0 49220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1490_
timestamp 1667941163
transform 1 0 48484 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1491_
timestamp 1667941163
transform 1 0 50324 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1492_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 52348 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1493_
timestamp 1667941163
transform -1 0 50324 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1494_
timestamp 1667941163
transform 1 0 50324 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1495_
timestamp 1667941163
transform -1 0 47656 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1496_
timestamp 1667941163
transform 1 0 40940 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1497_
timestamp 1667941163
transform -1 0 44712 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1498_
timestamp 1667941163
transform 1 0 49128 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1499_
timestamp 1667941163
transform 1 0 50784 0 -1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__o211a_1  _1500_
timestamp 1667941163
transform -1 0 46736 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1501_
timestamp 1667941163
transform 1 0 46644 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1502_
timestamp 1667941163
transform 1 0 48852 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1503_
timestamp 1667941163
transform 1 0 49312 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1504_
timestamp 1667941163
transform 1 0 50324 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1505_
timestamp 1667941163
transform 1 0 51428 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1506_
timestamp 1667941163
transform 1 0 52900 0 -1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1507_
timestamp 1667941163
transform -1 0 50416 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1508_
timestamp 1667941163
transform 1 0 50324 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1509_
timestamp 1667941163
transform 1 0 47748 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1510_
timestamp 1667941163
transform 1 0 50324 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__a2bb2o_1  _1511_
timestamp 1667941163
transform 1 0 52256 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1512_
timestamp 1667941163
transform 1 0 51796 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1513_
timestamp 1667941163
transform 1 0 51796 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1514_
timestamp 1667941163
transform 1 0 52992 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1515_
timestamp 1667941163
transform 1 0 53268 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1516_
timestamp 1667941163
transform -1 0 47840 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1517_
timestamp 1667941163
transform 1 0 48208 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1518_
timestamp 1667941163
transform 1 0 49036 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1519_
timestamp 1667941163
transform 1 0 50600 0 1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _1520_
timestamp 1667941163
transform 1 0 53360 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1521_
timestamp 1667941163
transform 1 0 54096 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1522_
timestamp 1667941163
transform 1 0 54556 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1523_
timestamp 1667941163
transform -1 0 56672 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__a22oi_1  _1524_
timestamp 1667941163
transform 1 0 51888 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1525_
timestamp 1667941163
transform 1 0 52900 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1526_
timestamp 1667941163
transform 1 0 52532 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1527_
timestamp 1667941163
transform 1 0 53728 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__a2bb2o_1  _1528_
timestamp 1667941163
transform 1 0 55476 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1529_
timestamp 1667941163
transform 1 0 54924 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1530_
timestamp 1667941163
transform -1 0 55016 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1531_
timestamp 1667941163
transform -1 0 54096 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1532_
timestamp 1667941163
transform 1 0 54096 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1533_
timestamp 1667941163
transform 1 0 53176 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1534_
timestamp 1667941163
transform 1 0 53912 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1535_
timestamp 1667941163
transform 1 0 52900 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1536_
timestamp 1667941163
transform 1 0 53176 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1537_
timestamp 1667941163
transform 1 0 54740 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1538_
timestamp 1667941163
transform -1 0 54740 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1539_
timestamp 1667941163
transform 1 0 55752 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1540_
timestamp 1667941163
transform -1 0 56580 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1541_
timestamp 1667941163
transform 1 0 55292 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1542_
timestamp 1667941163
transform -1 0 55936 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1543_
timestamp 1667941163
transform 1 0 55752 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1544_
timestamp 1667941163
transform -1 0 55384 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1545_
timestamp 1667941163
transform 1 0 53544 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1546_
timestamp 1667941163
transform -1 0 48944 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1547_
timestamp 1667941163
transform 1 0 48484 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1548_
timestamp 1667941163
transform -1 0 48944 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1549_
timestamp 1667941163
transform 1 0 47748 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1550_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 50968 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1551_
timestamp 1667941163
transform 1 0 50416 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1552_
timestamp 1667941163
transform 1 0 49128 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1553_
timestamp 1667941163
transform -1 0 50784 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1554_
timestamp 1667941163
transform -1 0 49864 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1555_
timestamp 1667941163
transform -1 0 51060 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1556_
timestamp 1667941163
transform -1 0 52256 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1557_
timestamp 1667941163
transform -1 0 51612 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1558_
timestamp 1667941163
transform 1 0 51888 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1559_
timestamp 1667941163
transform -1 0 51520 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1560_
timestamp 1667941163
transform 1 0 49772 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1561_
timestamp 1667941163
transform -1 0 48300 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1562_
timestamp 1667941163
transform -1 0 48300 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1563_
timestamp 1667941163
transform 1 0 47380 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1564_
timestamp 1667941163
transform -1 0 47932 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1565_
timestamp 1667941163
transform -1 0 47012 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1566_
timestamp 1667941163
transform -1 0 50600 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _1567_
timestamp 1667941163
transform 1 0 51152 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1568_
timestamp 1667941163
transform 1 0 50324 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1569_
timestamp 1667941163
transform 1 0 50876 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1570_
timestamp 1667941163
transform -1 0 51244 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1571_
timestamp 1667941163
transform 1 0 50324 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1572_
timestamp 1667941163
transform 1 0 47748 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1573_
timestamp 1667941163
transform 1 0 48760 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1574_
timestamp 1667941163
transform 1 0 48392 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1575_
timestamp 1667941163
transform -1 0 46460 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1576_
timestamp 1667941163
transform 1 0 46276 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1577_
timestamp 1667941163
transform 1 0 46092 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1578_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 44068 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1579_
timestamp 1667941163
transform -1 0 44620 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1580_
timestamp 1667941163
transform -1 0 45816 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1581_
timestamp 1667941163
transform -1 0 46828 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1582_
timestamp 1667941163
transform -1 0 46644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1583_
timestamp 1667941163
transform -1 0 46920 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1584_
timestamp 1667941163
transform -1 0 50508 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1585_
timestamp 1667941163
transform -1 0 50784 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1586_
timestamp 1667941163
transform 1 0 51152 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1587_
timestamp 1667941163
transform -1 0 36156 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1588_
timestamp 1667941163
transform -1 0 35972 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1589_
timestamp 1667941163
transform 1 0 40664 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1590_
timestamp 1667941163
transform -1 0 43516 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1591_
timestamp 1667941163
transform -1 0 37720 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1592_
timestamp 1667941163
transform 1 0 39100 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1593_
timestamp 1667941163
transform 1 0 45172 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1594_
timestamp 1667941163
transform 1 0 45172 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1595_
timestamp 1667941163
transform 1 0 51336 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1596_
timestamp 1667941163
transform -1 0 49312 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1597_
timestamp 1667941163
transform -1 0 49404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1598_
timestamp 1667941163
transform 1 0 47196 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1599_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 41676 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1600_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37904 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1601_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36432 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1602_
timestamp 1667941163
transform 1 0 40112 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1603_
timestamp 1667941163
transform 1 0 34868 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1604_
timestamp 1667941163
transform 1 0 38272 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1605_
timestamp 1667941163
transform -1 0 34224 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1606_
timestamp 1667941163
transform 1 0 31280 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1607_
timestamp 1667941163
transform 1 0 32292 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1608_
timestamp 1667941163
transform -1 0 33028 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1609_
timestamp 1667941163
transform -1 0 31648 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1610_
timestamp 1667941163
transform -1 0 30452 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1611_
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1612_
timestamp 1667941163
transform -1 0 30268 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1613_
timestamp 1667941163
transform -1 0 31924 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1614_
timestamp 1667941163
transform -1 0 42412 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1615_
timestamp 1667941163
transform 1 0 34868 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1616_
timestamp 1667941163
transform -1 0 31556 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1617_
timestamp 1667941163
transform -1 0 32660 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1618_
timestamp 1667941163
transform 1 0 29716 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1619_
timestamp 1667941163
transform 1 0 34592 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1620_
timestamp 1667941163
transform 1 0 32936 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1621_
timestamp 1667941163
transform 1 0 33396 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1622_
timestamp 1667941163
transform 1 0 33304 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1623_
timestamp 1667941163
transform 1 0 33120 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1624_
timestamp 1667941163
transform 1 0 41492 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1625_
timestamp 1667941163
transform 1 0 41952 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1626_
timestamp 1667941163
transform 1 0 43700 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1627_
timestamp 1667941163
transform -1 0 44252 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1628_
timestamp 1667941163
transform 1 0 43148 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1629_
timestamp 1667941163
transform 1 0 41124 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1630_
timestamp 1667941163
transform 1 0 44160 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_1  _1631_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 51244 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1632_ OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 50968 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_2  _1633_
timestamp 1667941163
transform 1 0 34776 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1634_
timestamp 1667941163
transform 1 0 34592 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1635_
timestamp 1667941163
transform 1 0 40020 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1636_
timestamp 1667941163
transform -1 0 42136 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1637_
timestamp 1667941163
transform 1 0 35972 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1638_
timestamp 1667941163
transform 1 0 38088 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1639_
timestamp 1667941163
transform 1 0 43976 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1640_
timestamp 1667941163
transform 1 0 43792 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1641_
timestamp 1667941163
transform -1 0 51888 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1642_
timestamp 1667941163
transform 1 0 47380 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1643_
timestamp 1667941163
transform 1 0 48024 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1644_
timestamp 1667941163
transform 1 0 46184 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_net8 OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34776 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_net12
timestamp 1667941163
transform 1 0 48760 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_net8
timestamp 1667941163
transform -1 0 33028 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_net12
timestamp 1667941163
transform -1 0 48668 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_net8
timestamp 1667941163
transform -1 0 33856 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_net12
timestamp 1667941163
transform 1 0 50324 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout8
timestamp 1667941163
transform 1 0 29900 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout9
timestamp 1667941163
transform 1 0 28060 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout10
timestamp 1667941163
transform 1 0 27324 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout11
timestamp 1667941163
transform -1 0 43516 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout12
timestamp 1667941163
transform 1 0 47748 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout13
timestamp 1667941163
transform 1 0 40756 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 OSPDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 39100 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1667941163
transform -1 0 58420 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform -1 0 1840 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1667941163
transform -1 0 58420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1667941163
transform 1 0 58052 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1667941163
transform -1 0 1932 0 1 30464
box -38 -48 406 592
<< labels >>
flabel metal2 s 59910 59200 59966 59800 0 FreeSans 224 90 0 0 A_PAD
port 0 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 B_PAD
port 1 nsew signal input
flabel metal3 s 59200 29248 59800 29368 0 FreeSans 480 0 0 0 OUT_1
port 2 nsew signal tristate
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 OUT_2
port 3 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 sel
port 4 nsew signal input
flabel metal2 s 1306 59200 1362 59800 0 FreeSans 224 90 0 0 user_clock2
port 5 nsew signal input
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 6 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 6 nsew power bidirectional
flabel metal5 s 1056 5346 58928 5666 0 FreeSans 2560 0 0 0 vccd1
port 6 nsew power bidirectional
flabel metal5 s 1056 35982 58928 36302 0 FreeSans 2560 0 0 0 vccd1
port 6 nsew power bidirectional
flabel metal4 s 4868 2128 5188 57712 0 FreeSans 1920 90 0 0 vssd1
port 7 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 57712 0 FreeSans 1920 90 0 0 vssd1
port 7 nsew ground bidirectional
flabel metal5 s 1056 6006 58928 6326 0 FreeSans 2560 0 0 0 vssd1
port 7 nsew ground bidirectional
flabel metal5 s 1056 36642 58928 36962 0 FreeSans 2560 0 0 0 vssd1
port 7 nsew ground bidirectional
flabel metal2 s 30930 59200 30986 59800 0 FreeSans 224 90 0 0 wb_clk_i
port 8 nsew signal input
flabel metal2 s 58622 200 58678 800 0 FreeSans 224 90 0 0 wb_rst_i
port 9 nsew signal input
rlabel metal1 29992 57120 29992 57120 0 vccd1
rlabel metal1 29992 57664 29992 57664 0 vssd1
rlabel metal1 59110 56814 59110 56814 0 A_PAD
rlabel metal1 29072 2278 29072 2278 0 B_PAD
rlabel metal1 43378 27642 43378 27642 0 MUL.PS_R1_inst1.LUT_inst1.i0
rlabel metal1 38824 33898 38824 33898 0 MUL.PS_R1_inst1.LUT_inst1.i1
rlabel metal2 36662 26962 36662 26962 0 MUL.PS_R1_inst1.LUT_inst1.i3
rlabel metal2 30682 34612 30682 34612 0 MUL.PS_R1_inst1.LUT_inst1.i4
rlabel metal1 31188 31994 31188 31994 0 MUL.PS_R1_inst1.LUT_inst10.I0
rlabel metal1 29624 29818 29624 29818 0 MUL.PS_R1_inst1.LUT_inst10.I1
rlabel metal1 28704 36006 28704 36006 0 MUL.PS_R1_inst1.LUT_inst11.I1
rlabel metal2 30222 36210 30222 36210 0 MUL.PS_R1_inst1.LUT_inst12.I1
rlabel metal1 28382 31450 28382 31450 0 MUL.PS_R1_inst1.LUT_inst13.I1
rlabel metal1 29670 30770 29670 30770 0 MUL.PS_R1_inst1.LUT_inst14.I1
rlabel metal1 40296 34034 40296 34034 0 MUL.PS_R1_inst1.LUT_inst15.I1
rlabel metal1 38824 30838 38824 30838 0 MUL.PS_R1_inst1.LUT_inst2.I1
rlabel via2 41906 33099 41906 33099 0 MUL.PS_R1_inst1.LUT_inst3.I1
rlabel metal1 37030 34170 37030 34170 0 MUL.PS_R1_inst1.LUT_inst4.I1
rlabel metal1 37306 48042 37306 48042 0 MUL.PS_R1_inst1.LUT_inst5.I1
rlabel metal2 32430 30141 32430 30141 0 MUL.PS_R1_inst1.LUT_inst6.I1
rlabel metal1 33626 33082 33626 33082 0 MUL.PS_R1_inst1.LUT_inst7.I1
rlabel metal1 31326 46002 31326 46002 0 MUL.PS_R1_inst1.LUT_inst8.I1
rlabel metal1 33166 35054 33166 35054 0 MUL.PS_Rx_inst2.LUT_inst1.i3
rlabel metal2 32890 36210 32890 36210 0 MUL.PS_Rx_inst2.LUT_inst1.i4
rlabel metal1 35834 30634 35834 30634 0 MUL.PS_Rx_inst3.LUT_inst1.i3
rlabel metal2 34730 33014 34730 33014 0 MUL.PS_Rx_inst3.LUT_inst1.i4
rlabel via1 35558 34595 35558 34595 0 MUL.PS_Rx_inst4.LUT_inst1.i3
rlabel metal1 35512 32402 35512 32402 0 MUL.PS_Rx_inst4.LUT_inst1.i4
rlabel metal1 36892 26962 36892 26962 0 MUL.PS_Rx_inst5.LUT_inst1.i3
rlabel metal1 43608 36142 43608 36142 0 MUL.PS_Rx_inst5.LUT_inst1.i4
rlabel via2 44022 29597 44022 29597 0 MUL.PS_Rx_inst6.LUT_inst1.i3
rlabel metal2 46046 32912 46046 32912 0 MUL.PS_Rx_inst6.LUT_inst1.i4
rlabel metal1 46506 34510 46506 34510 0 MUL.PS_Rx_inst7.LUT_inst1.i3
rlabel metal1 48438 33830 48438 33830 0 MUL.PS_Rx_inst7.LUT_inst1.i4
rlabel metal1 41722 28492 41722 28492 0 MUL.PS_Rx_inst8.LUT_inst1.i3
rlabel metal1 47840 31858 47840 31858 0 MUL.PS_Rx_inst8.LUT_inst1.i4
rlabel metal2 58282 29393 58282 29393 0 OUT_1
rlabel metal3 1188 30668 1188 30668 0 OUT_2
rlabel metal1 42872 27846 42872 27846 0 _0000_
rlabel metal1 39008 33082 39008 33082 0 _0001_
rlabel metal1 37536 31110 37536 31110 0 _0002_
rlabel metal2 41446 33048 41446 33048 0 _0003_
rlabel metal2 36202 34136 36202 34136 0 _0004_
rlabel metal1 39376 34170 39376 34170 0 _0005_
rlabel metal1 32752 29274 32752 29274 0 _0006_
rlabel metal1 33265 32810 33265 32810 0 _0007_
rlabel metal2 33166 28254 33166 28254 0 _0008_
rlabel metal2 32430 31586 32430 31586 0 _0009_
rlabel metal2 30222 29444 30222 29444 0 _0010_
rlabel metal2 29670 32606 29670 32606 0 _0011_
rlabel metal2 29118 34408 29118 34408 0 _0012_
rlabel metal1 29677 31382 29677 31382 0 _0013_
rlabel metal2 30866 30464 30866 30464 0 _0014_
rlabel metal2 41998 33762 41998 33762 0 _0015_
rlabel metal1 35880 25466 35880 25466 0 _0016_
rlabel metal2 30590 33490 30590 33490 0 _0017_
rlabel metal2 31694 28696 31694 28696 0 _0018_
rlabel metal1 31004 32538 31004 32538 0 _0019_
rlabel metal1 35190 29818 35190 29818 0 _0020_
rlabel metal1 34224 31994 34224 31994 0 _0021_
rlabel metal1 34914 28730 34914 28730 0 _0022_
rlabel metal1 34086 31858 34086 31858 0 _0023_
rlabel metal1 34224 26554 34224 26554 0 _0024_
rlabel metal1 43247 30634 43247 30634 0 _0025_
rlabel metal1 43424 29274 43424 29274 0 _0026_
rlabel metal2 44482 32606 44482 32606 0 _0027_
rlabel metal2 43654 26146 43654 26146 0 _0028_
rlabel metal2 44574 30022 44574 30022 0 _0029_
rlabel metal1 43286 24378 43286 24378 0 _0030_
rlabel metal1 44843 22678 44843 22678 0 _0031_
rlabel metal1 36064 23222 36064 23222 0 _0032_
rlabel metal1 35926 24378 35926 24378 0 _0033_
rlabel metal2 40802 22882 40802 22882 0 _0034_
rlabel metal1 43056 23562 43056 23562 0 _0035_
rlabel metal2 37582 21794 37582 21794 0 _0036_
rlabel metal1 39192 21658 39192 21658 0 _0037_
rlabel metal2 45310 23902 45310 23902 0 _0038_
rlabel metal1 45264 25126 45264 25126 0 _0039_
rlabel metal1 51297 23766 51297 23766 0 _0040_
rlabel metal1 49128 23834 49128 23834 0 _0041_
rlabel metal1 49358 22066 49358 22066 0 _0042_
rlabel metal1 47242 22066 47242 22066 0 _0043_
rlabel metal1 42083 27642 42083 27642 0 _0044_
rlabel metal1 38134 32538 38134 32538 0 _0045_
rlabel metal2 36478 30192 36478 30192 0 _0046_
rlabel metal1 40618 32538 40618 32538 0 _0047_
rlabel metal2 36570 33558 36570 33558 0 _0048_
rlabel metal2 39146 33456 39146 33456 0 _0049_
rlabel metal1 34316 30294 34316 30294 0 _0050_
rlabel metal2 31602 32674 31602 32674 0 _0051_
rlabel metal2 32614 27812 32614 27812 0 _0052_
rlabel metal1 38180 31246 38180 31246 0 _0053_
rlabel metal1 39330 29240 39330 29240 0 _0054_
rlabel metal1 34086 31960 34086 31960 0 _0055_
rlabel metal1 28612 30090 28612 30090 0 _0056_
rlabel metal1 37996 30770 37996 30770 0 _0057_
rlabel metal2 31694 30124 31694 30124 0 _0058_
rlabel metal2 41722 34476 41722 34476 0 _0059_
rlabel metal2 35190 26146 35190 26146 0 _0060_
rlabel metal1 36478 31994 36478 31994 0 _0061_
rlabel metal1 33074 28458 33074 28458 0 _0062_
rlabel metal1 36984 33014 36984 33014 0 _0063_
rlabel metal1 34914 30328 34914 30328 0 _0064_
rlabel metal1 34776 32334 34776 32334 0 _0065_
rlabel metal1 34730 28594 34730 28594 0 _0066_
rlabel metal2 33718 31076 33718 31076 0 _0067_
rlabel metal2 33442 27166 33442 27166 0 _0068_
rlabel metal2 41814 30872 41814 30872 0 _0069_
rlabel metal2 41722 29410 41722 29410 0 _0070_
rlabel metal1 42918 32470 42918 32470 0 _0071_
rlabel metal2 43930 26792 43930 26792 0 _0072_
rlabel metal1 42596 30158 42596 30158 0 _0073_
rlabel metal2 41078 26792 41078 26792 0 _0074_
rlabel metal2 44482 22814 44482 22814 0 _0075_
rlabel metal2 51106 24956 51106 24956 0 _0076_
rlabel via1 51285 26350 51285 26350 0 _0077_
rlabel metal2 35098 23902 35098 23902 0 _0078_
rlabel metal1 36202 24718 36202 24718 0 _0079_
rlabel metal1 38916 22066 38916 22066 0 _0080_
rlabel metal1 42228 23630 42228 23630 0 _0081_
rlabel via1 36287 22202 36287 22202 0 _0082_
rlabel metal1 38364 21658 38364 21658 0 _0083_
rlabel metal1 44298 23800 44298 23800 0 _0084_
rlabel metal1 44160 24718 44160 24718 0 _0085_
rlabel metal1 49634 23222 49634 23222 0 _0086_
rlabel metal2 47702 25262 47702 25262 0 _0087_
rlabel metal1 48438 22202 48438 22202 0 _0088_
rlabel metal1 46598 22746 46598 22746 0 _0089_
rlabel metal2 46874 23052 46874 23052 0 _0090_
rlabel metal1 48392 21998 48392 21998 0 _0091_
rlabel metal1 47242 26928 47242 26928 0 _0092_
rlabel metal2 49450 29036 49450 29036 0 _0093_
rlabel metal1 46000 26962 46000 26962 0 _0094_
rlabel metal1 37950 23698 37950 23698 0 _0095_
rlabel metal2 40066 25296 40066 25296 0 _0096_
rlabel metal1 46966 24650 46966 24650 0 _0097_
rlabel metal1 49726 25942 49726 25942 0 _0098_
rlabel metal2 48898 24412 48898 24412 0 _0099_
rlabel metal1 48208 25874 48208 25874 0 _0100_
rlabel via1 45696 28526 45696 28526 0 _0101_
rlabel metal2 56258 35292 56258 35292 0 _0102_
rlabel metal1 45172 25874 45172 25874 0 _0103_
rlabel metal2 51658 34918 51658 34918 0 _0104_
rlabel metal1 53084 33490 53084 33490 0 _0105_
rlabel metal2 46322 24684 46322 24684 0 _0106_
rlabel metal1 38548 22950 38548 22950 0 _0107_
rlabel metal1 38410 21522 38410 21522 0 _0108_
rlabel metal1 36432 22610 36432 22610 0 _0109_
rlabel metal2 39054 24922 39054 24922 0 _0110_
rlabel metal1 36938 25194 36938 25194 0 _0111_
rlabel metal1 40756 26418 40756 26418 0 _0112_
rlabel metal1 39606 24582 39606 24582 0 _0113_
rlabel metal2 39146 25738 39146 25738 0 _0114_
rlabel metal2 38042 25636 38042 25636 0 _0115_
rlabel metal2 40066 28832 40066 28832 0 _0116_
rlabel metal1 38410 25908 38410 25908 0 _0117_
rlabel metal1 38732 25670 38732 25670 0 _0118_
rlabel metal1 38732 21998 38732 21998 0 _0119_
rlabel metal1 42826 23732 42826 23732 0 _0120_
rlabel metal1 37904 23834 37904 23834 0 _0121_
rlabel metal1 39284 23766 39284 23766 0 _0122_
rlabel metal1 38318 23494 38318 23494 0 _0123_
rlabel metal2 38870 23562 38870 23562 0 _0124_
rlabel metal1 35282 24208 35282 24208 0 _0125_
rlabel metal1 45034 23086 45034 23086 0 _0126_
rlabel viali 39874 24854 39874 24854 0 _0127_
rlabel metal1 41285 27438 41285 27438 0 _0128_
rlabel metal1 40940 27642 40940 27642 0 _0129_
rlabel metal1 37766 29546 37766 29546 0 _0130_
rlabel metal1 41216 28526 41216 28526 0 _0131_
rlabel metal2 42734 28764 42734 28764 0 _0132_
rlabel metal1 38548 28390 38548 28390 0 _0133_
rlabel metal1 36846 31824 36846 31824 0 _0134_
rlabel via1 40539 30634 40539 30634 0 _0135_
rlabel metal1 48668 31790 48668 31790 0 _0136_
rlabel metal1 39836 26962 39836 26962 0 _0137_
rlabel metal1 39514 26996 39514 26996 0 _0138_
rlabel metal2 41354 27506 41354 27506 0 _0139_
rlabel metal1 43010 26554 43010 26554 0 _0140_
rlabel metal1 46046 33286 46046 33286 0 _0141_
rlabel metal2 40250 31994 40250 31994 0 _0142_
rlabel metal1 38824 31110 38824 31110 0 _0143_
rlabel metal2 38870 32096 38870 32096 0 _0144_
rlabel metal1 38686 32946 38686 32946 0 _0145_
rlabel metal2 37306 27744 37306 27744 0 _0146_
rlabel metal1 40250 28186 40250 28186 0 _0147_
rlabel metal2 39054 27472 39054 27472 0 _0148_
rlabel metal1 40549 31382 40549 31382 0 _0149_
rlabel metal1 43102 33830 43102 33830 0 _0150_
rlabel metal2 36294 26452 36294 26452 0 _0151_
rlabel metal1 34730 27098 34730 27098 0 _0152_
rlabel metal2 38962 37366 38962 37366 0 _0153_
rlabel metal1 33948 30702 33948 30702 0 _0154_
rlabel metal2 39698 25500 39698 25500 0 _0155_
rlabel metal2 39238 26894 39238 26894 0 _0156_
rlabel metal1 39836 32470 39836 32470 0 _0157_
rlabel metal1 38870 28424 38870 28424 0 _0158_
rlabel metal1 39560 27574 39560 27574 0 _0159_
rlabel metal1 34592 33286 34592 33286 0 _0160_
rlabel metal1 35558 27030 35558 27030 0 _0161_
rlabel metal1 33074 30668 33074 30668 0 _0162_
rlabel metal1 38180 32810 38180 32810 0 _0163_
rlabel metal2 33810 33762 33810 33762 0 _0164_
rlabel metal1 36892 28730 36892 28730 0 _0165_
rlabel metal1 37191 31722 37191 31722 0 _0166_
rlabel metal2 37214 32334 37214 32334 0 _0167_
rlabel metal1 35420 25874 35420 25874 0 _0168_
rlabel via1 36845 38930 36845 38930 0 _0169_
rlabel metal1 41860 34578 41860 34578 0 _0170_
rlabel metal2 41170 34782 41170 34782 0 _0171_
rlabel metal2 39974 29682 39974 29682 0 _0172_
rlabel metal1 40112 36142 40112 36142 0 _0173_
rlabel metal1 51520 32878 51520 32878 0 _0174_
rlabel metal1 40020 30702 40020 30702 0 _0175_
rlabel metal1 32522 38250 32522 38250 0 _0176_
rlabel metal1 40710 37638 40710 37638 0 _0177_
rlabel metal1 38686 40018 38686 40018 0 _0178_
rlabel metal1 51934 36856 51934 36856 0 _0179_
rlabel metal2 28842 29852 28842 29852 0 _0180_
rlabel metal2 35558 40868 35558 40868 0 _0181_
rlabel metal1 54832 35666 54832 35666 0 _0182_
rlabel metal2 40434 32096 40434 32096 0 _0183_
rlabel metal1 39836 41106 39836 41106 0 _0184_
rlabel metal1 40664 40358 40664 40358 0 _0185_
rlabel metal1 31234 45424 31234 45424 0 _0186_
rlabel metal1 40618 31212 40618 31212 0 _0187_
rlabel metal1 40986 44302 40986 44302 0 _0188_
rlabel metal2 36570 35564 36570 35564 0 _0189_
rlabel metal1 32798 27472 32798 27472 0 _0190_
rlabel metal1 36708 43690 36708 43690 0 _0191_
rlabel metal1 36087 31790 36087 31790 0 _0192_
rlabel metal2 35374 32096 35374 32096 0 _0193_
rlabel metal2 41354 43826 41354 43826 0 _0194_
rlabel metal2 38180 36516 38180 36516 0 _0195_
rlabel metal1 40802 45832 40802 45832 0 _0196_
rlabel metal1 41216 31994 41216 31994 0 _0197_
rlabel metal2 38870 45220 38870 45220 0 _0198_
rlabel via2 37582 32555 37582 32555 0 _0199_
rlabel metal1 36432 32878 36432 32878 0 _0200_
rlabel metal2 38226 44608 38226 44608 0 _0201_
rlabel metal2 37582 41004 37582 41004 0 _0202_
rlabel metal1 48438 41106 48438 41106 0 _0203_
rlabel metal2 37582 35343 37582 35343 0 _0204_
rlabel metal1 53590 32402 53590 32402 0 _0205_
rlabel metal2 44942 25024 44942 25024 0 _0206_
rlabel metal2 41814 28356 41814 28356 0 _0207_
rlabel metal1 1656 56406 1656 56406 0 _0208_
rlabel metal1 47150 21998 47150 21998 0 _0209_
rlabel metal1 33718 32538 33718 32538 0 _0210_
rlabel metal1 30498 29138 30498 29138 0 _0211_
rlabel metal1 34500 31790 34500 31790 0 _0212_
rlabel metal1 39146 21488 39146 21488 0 _0213_
rlabel metal1 51566 24718 51566 24718 0 _0214_
rlabel metal2 35374 35122 35374 35122 0 _0215_
rlabel metal1 37122 37774 37122 37774 0 _0216_
rlabel via1 35463 41106 35463 41106 0 _0217_
rlabel via1 40963 38318 40963 38318 0 _0218_
rlabel metal1 35282 39338 35282 39338 0 _0219_
rlabel metal1 41354 39542 41354 39542 0 _0220_
rlabel metal1 34960 40698 34960 40698 0 _0221_
rlabel metal1 36846 40698 36846 40698 0 _0222_
rlabel metal1 35512 38862 35512 38862 0 _0223_
rlabel metal1 37168 40562 37168 40562 0 _0224_
rlabel metal1 39744 43282 39744 43282 0 _0225_
rlabel metal2 40618 43588 40618 43588 0 _0226_
rlabel metal1 40434 37400 40434 37400 0 _0227_
rlabel metal1 33028 36550 33028 36550 0 _0228_
rlabel metal1 35098 36890 35098 36890 0 _0229_
rlabel metal1 32844 38930 32844 38930 0 _0230_
rlabel via1 38755 41106 38755 41106 0 _0231_
rlabel metal1 31050 40120 31050 40120 0 _0232_
rlabel metal1 32936 37978 32936 37978 0 _0233_
rlabel metal2 32338 38386 32338 38386 0 _0234_
rlabel metal2 37030 40052 37030 40052 0 _0235_
rlabel metal2 32798 38216 32798 38216 0 _0236_
rlabel metal2 37858 40018 37858 40018 0 _0237_
rlabel metal2 38594 46716 38594 46716 0 _0238_
rlabel metal1 39100 46682 39100 46682 0 _0239_
rlabel metal2 31234 36754 31234 36754 0 _0240_
rlabel metal1 33534 35802 33534 35802 0 _0241_
rlabel metal1 31901 36142 31901 36142 0 _0242_
rlabel metal2 32844 41400 32844 41400 0 _0243_
rlabel metal1 32844 34510 32844 34510 0 _0244_
rlabel metal1 29670 35258 29670 35258 0 _0245_
rlabel metal1 31878 41582 31878 41582 0 _0246_
rlabel metal1 34178 37366 34178 37366 0 _0247_
rlabel metal1 31464 45458 31464 45458 0 _0248_
rlabel metal2 32798 35972 32798 35972 0 _0249_
rlabel metal1 30820 45458 30820 45458 0 _0250_
rlabel metal1 34684 45322 34684 45322 0 _0251_
rlabel metal2 36018 47056 36018 47056 0 _0252_
rlabel metal1 37260 45322 37260 45322 0 _0253_
rlabel metal2 37766 46784 37766 46784 0 _0254_
rlabel metal1 38042 47532 38042 47532 0 _0255_
rlabel metal2 40158 46274 40158 46274 0 _0256_
rlabel metal1 38180 43758 38180 43758 0 _0257_
rlabel metal1 38962 43656 38962 43656 0 _0258_
rlabel metal2 36938 44540 36938 44540 0 _0259_
rlabel metal2 37858 43758 37858 43758 0 _0260_
rlabel metal2 38962 44812 38962 44812 0 _0261_
rlabel metal1 40572 35666 40572 35666 0 _0262_
rlabel metal2 40710 43996 40710 43996 0 _0263_
rlabel metal3 41055 42908 41055 42908 0 _0264_
rlabel metal1 40112 45458 40112 45458 0 _0265_
rlabel metal2 40986 47022 40986 47022 0 _0266_
rlabel metal2 37490 46750 37490 46750 0 _0267_
rlabel metal1 37904 46682 37904 46682 0 _0268_
rlabel metal2 34638 46342 34638 46342 0 _0269_
rlabel metal1 33902 48110 33902 48110 0 _0270_
rlabel metal1 37030 48246 37030 48246 0 _0271_
rlabel metal2 38778 48382 38778 48382 0 _0272_
rlabel metal2 40618 48484 40618 48484 0 _0273_
rlabel metal2 43332 37196 43332 37196 0 _0274_
rlabel metal1 43056 35666 43056 35666 0 _0275_
rlabel metal1 41492 35802 41492 35802 0 _0276_
rlabel metal2 42918 38420 42918 38420 0 _0277_
rlabel metal1 43562 36550 43562 36550 0 _0278_
rlabel metal1 42734 34918 42734 34918 0 _0279_
rlabel metal2 43286 34646 43286 34646 0 _0280_
rlabel metal1 43516 34986 43516 34986 0 _0281_
rlabel metal2 43562 34850 43562 34850 0 _0282_
rlabel metal2 44206 34204 44206 34204 0 _0283_
rlabel metal1 45126 34102 45126 34102 0 _0284_
rlabel metal2 47242 30498 47242 30498 0 _0285_
rlabel via1 43104 37842 43104 37842 0 _0286_
rlabel metal1 44229 45934 44229 45934 0 _0287_
rlabel metal2 41538 36788 41538 36788 0 _0288_
rlabel metal1 43930 40426 43930 40426 0 _0289_
rlabel metal1 42458 37264 42458 37264 0 _0290_
rlabel metal1 42044 40494 42044 40494 0 _0291_
rlabel metal1 43562 45594 43562 45594 0 _0292_
rlabel metal1 44390 46138 44390 46138 0 _0293_
rlabel metal2 40434 46410 40434 46410 0 _0294_
rlabel metal1 41170 46138 41170 46138 0 _0295_
rlabel metal2 31142 45050 31142 45050 0 _0296_
rlabel metal1 31464 44370 31464 44370 0 _0297_
rlabel metal2 32338 46410 32338 46410 0 _0298_
rlabel metal1 32752 46138 32752 46138 0 _0299_
rlabel metal2 31786 46342 31786 46342 0 _0300_
rlabel metal2 32614 47838 32614 47838 0 _0301_
rlabel metal1 33166 47566 33166 47566 0 _0302_
rlabel metal1 35742 47532 35742 47532 0 _0303_
rlabel metal1 34914 46988 34914 46988 0 _0304_
rlabel metal1 35604 46886 35604 46886 0 _0305_
rlabel metal1 34592 48178 34592 48178 0 _0306_
rlabel metal1 36294 48722 36294 48722 0 _0307_
rlabel metal1 40710 48178 40710 48178 0 _0308_
rlabel metal2 42918 48144 42918 48144 0 _0309_
rlabel metal1 39468 46546 39468 46546 0 _0310_
rlabel metal1 40296 46682 40296 46682 0 _0311_
rlabel metal1 39054 48620 39054 48620 0 _0312_
rlabel metal1 42918 48620 42918 48620 0 _0313_
rlabel metal2 44298 48076 44298 48076 0 _0314_
rlabel metal1 45954 34578 45954 34578 0 _0315_
rlabel metal1 46828 36142 46828 36142 0 _0316_
rlabel metal2 46506 36890 46506 36890 0 _0317_
rlabel metal2 48162 35530 48162 35530 0 _0318_
rlabel via1 48532 39406 48532 39406 0 _0319_
rlabel metal1 49082 36822 49082 36822 0 _0320_
rlabel metal1 45034 36142 45034 36142 0 _0321_
rlabel metal1 45586 35802 45586 35802 0 _0322_
rlabel metal2 45218 36380 45218 36380 0 _0323_
rlabel metal2 45126 35530 45126 35530 0 _0324_
rlabel metal1 45678 34442 45678 34442 0 _0325_
rlabel metal1 46506 29138 46506 29138 0 _0326_
rlabel metal2 44206 42874 44206 42874 0 _0327_
rlabel metal1 44712 43282 44712 43282 0 _0328_
rlabel metal2 44390 45866 44390 45866 0 _0329_
rlabel via2 46966 31331 46966 31331 0 _0330_
rlabel metal2 46966 30124 46966 30124 0 _0331_
rlabel metal1 52992 28458 52992 28458 0 _0332_
rlabel metal1 46782 28934 46782 28934 0 _0333_
rlabel metal1 49450 26316 49450 26316 0 _0334_
rlabel metal2 32890 44676 32890 44676 0 _0335_
rlabel metal1 33948 44370 33948 44370 0 _0336_
rlabel metal1 30958 41616 30958 41616 0 _0337_
rlabel metal1 30912 43282 30912 43282 0 _0338_
rlabel metal1 33534 44268 33534 44268 0 _0339_
rlabel metal1 35742 44846 35742 44846 0 _0340_
rlabel metal1 35098 42636 35098 42636 0 _0341_
rlabel metal1 35650 42534 35650 42534 0 _0342_
rlabel metal2 31786 42500 31786 42500 0 _0343_
rlabel metal2 32706 43282 32706 43282 0 _0344_
rlabel metal2 29946 36550 29946 36550 0 _0345_
rlabel metal1 29946 42194 29946 42194 0 _0346_
rlabel metal2 31142 43486 31142 43486 0 _0347_
rlabel metal1 35190 44336 35190 44336 0 _0348_
rlabel metal2 35374 45084 35374 45084 0 _0349_
rlabel metal2 45034 45118 45034 45118 0 _0350_
rlabel metal2 42090 45934 42090 45934 0 _0351_
rlabel metal2 43286 46852 43286 46852 0 _0352_
rlabel metal1 40572 46546 40572 46546 0 _0353_
rlabel metal1 40986 47600 40986 47600 0 _0354_
rlabel metal1 37076 47498 37076 47498 0 _0355_
rlabel metal1 41354 47702 41354 47702 0 _0356_
rlabel metal2 45034 46852 45034 46852 0 _0357_
rlabel metal1 48070 46580 48070 46580 0 _0358_
rlabel metal2 42642 43452 42642 43452 0 _0359_
rlabel metal1 43378 43418 43378 43418 0 _0360_
rlabel metal1 34868 42330 34868 42330 0 _0361_
rlabel metal2 33994 43180 33994 43180 0 _0362_
rlabel metal1 30774 40052 30774 40052 0 _0363_
rlabel metal1 31142 42670 31142 42670 0 _0364_
rlabel metal2 29210 37230 29210 37230 0 _0365_
rlabel metal1 29072 41582 29072 41582 0 _0366_
rlabel metal2 30222 42432 30222 42432 0 _0367_
rlabel metal2 32982 43078 32982 43078 0 _0368_
rlabel metal1 34454 43418 34454 43418 0 _0369_
rlabel metal1 43654 44404 43654 44404 0 _0370_
rlabel metal2 43838 45220 43838 45220 0 _0371_
rlabel metal1 47978 45390 47978 45390 0 _0372_
rlabel metal1 48484 37162 48484 37162 0 _0373_
rlabel metal1 53314 38862 53314 38862 0 _0374_
rlabel metal2 46966 37638 46966 37638 0 _0375_
rlabel metal1 49542 38930 49542 38930 0 _0376_
rlabel metal2 47794 36992 47794 36992 0 _0377_
rlabel metal2 51658 39168 51658 39168 0 _0378_
rlabel metal1 47794 44302 47794 44302 0 _0379_
rlabel metal2 48438 44948 48438 44948 0 _0380_
rlabel metal1 48438 45594 48438 45594 0 _0381_
rlabel metal1 49634 40052 49634 40052 0 _0382_
rlabel metal1 48622 43146 48622 43146 0 _0383_
rlabel metal2 49266 43962 49266 43962 0 _0384_
rlabel metal1 36984 42874 36984 42874 0 _0385_
rlabel metal1 37030 43418 37030 43418 0 _0386_
rlabel metal1 29854 39542 29854 39542 0 _0387_
rlabel metal1 30498 41582 30498 41582 0 _0388_
rlabel metal1 29440 37230 29440 37230 0 _0389_
rlabel metal1 28888 40494 28888 40494 0 _0390_
rlabel metal1 29624 41650 29624 41650 0 _0391_
rlabel metal1 30498 41480 30498 41480 0 _0392_
rlabel metal1 35512 43146 35512 43146 0 _0393_
rlabel via2 45402 43741 45402 43741 0 _0394_
rlabel metal2 41998 43452 41998 43452 0 _0395_
rlabel metal1 43194 43962 43194 43962 0 _0396_
rlabel metal2 44022 44574 44022 44574 0 _0397_
rlabel metal1 48990 44914 48990 44914 0 _0398_
rlabel metal2 49174 44268 49174 44268 0 _0399_
rlabel metal1 50324 43282 50324 43282 0 _0400_
rlabel metal1 53774 35020 53774 35020 0 _0401_
rlabel metal1 52118 39950 52118 39950 0 _0402_
rlabel metal2 48714 34272 48714 34272 0 _0403_
rlabel metal1 48530 33898 48530 33898 0 _0404_
rlabel metal1 54970 35734 54970 35734 0 _0405_
rlabel metal2 52118 35462 52118 35462 0 _0406_
rlabel metal2 49266 41990 49266 41990 0 _0407_
rlabel metal1 53590 35156 53590 35156 0 _0408_
rlabel metal1 53590 36686 53590 36686 0 _0409_
rlabel metal1 50094 41650 50094 41650 0 _0410_
rlabel metal2 50922 41004 50922 41004 0 _0411_
rlabel metal1 51612 34578 51612 34578 0 _0412_
rlabel metal1 51014 30736 51014 30736 0 _0413_
rlabel metal2 51198 30532 51198 30532 0 _0414_
rlabel metal2 54326 32309 54326 32309 0 _0415_
rlabel metal1 55706 32844 55706 32844 0 _0416_
rlabel via1 49082 31994 49082 31994 0 _0417_
rlabel metal1 48806 30804 48806 30804 0 _0418_
rlabel metal2 51566 31110 51566 31110 0 _0419_
rlabel metal2 51382 30124 51382 30124 0 _0420_
rlabel metal1 51474 29070 51474 29070 0 _0421_
rlabel metal1 51382 28526 51382 28526 0 _0422_
rlabel metal1 45770 34034 45770 34034 0 _0423_
rlabel metal1 54418 37128 54418 37128 0 _0424_
rlabel metal2 48990 40698 48990 40698 0 _0425_
rlabel metal1 48622 40052 48622 40052 0 _0426_
rlabel metal1 47334 43418 47334 43418 0 _0427_
rlabel metal1 46690 43962 46690 43962 0 _0428_
rlabel metal2 43930 45407 43930 45407 0 _0429_
rlabel metal1 44942 46682 44942 46682 0 _0430_
rlabel metal1 44206 47090 44206 47090 0 _0431_
rlabel metal1 46414 47090 46414 47090 0 _0432_
rlabel metal2 47886 46988 47886 46988 0 _0433_
rlabel metal1 48438 39950 48438 39950 0 _0434_
rlabel metal1 48990 39916 48990 39916 0 _0435_
rlabel metal1 50094 39882 50094 39882 0 _0436_
rlabel metal2 47426 44370 47426 44370 0 _0437_
rlabel metal1 48438 42160 48438 42160 0 _0438_
rlabel metal2 47518 41820 47518 41820 0 _0439_
rlabel metal2 48024 38692 48024 38692 0 _0440_
rlabel metal1 50048 28730 50048 28730 0 _0441_
rlabel metal2 49174 28764 49174 28764 0 _0442_
rlabel metal2 47886 33864 47886 33864 0 _0443_
rlabel metal1 45724 33354 45724 33354 0 _0444_
rlabel metal1 46368 33966 46368 33966 0 _0445_
rlabel metal2 46230 33388 46230 33388 0 _0446_
rlabel metal1 47334 32980 47334 32980 0 _0447_
rlabel metal1 48024 29614 48024 29614 0 _0448_
rlabel metal1 46460 27302 46460 27302 0 _0449_
rlabel metal2 49082 29138 49082 29138 0 _0450_
rlabel metal2 49358 27370 49358 27370 0 _0451_
rlabel metal2 51198 25534 51198 25534 0 _0452_
rlabel metal2 35466 35394 35466 35394 0 _0453_
rlabel metal1 37076 35734 37076 35734 0 _0454_
rlabel metal1 38318 35564 38318 35564 0 _0455_
rlabel metal1 39606 35564 39606 35564 0 _0456_
rlabel metal1 40802 35530 40802 35530 0 _0457_
rlabel metal2 37950 40902 37950 40902 0 _0458_
rlabel metal1 38916 41242 38916 41242 0 _0459_
rlabel metal1 37628 41582 37628 41582 0 _0460_
rlabel metal2 38042 39043 38042 39043 0 _0461_
rlabel metal2 38870 42466 38870 42466 0 _0462_
rlabel via2 46966 26027 46966 26027 0 _0463_
rlabel metal1 44758 28118 44758 28118 0 _0464_
rlabel metal1 34592 36346 34592 36346 0 _0465_
rlabel metal1 35144 36618 35144 36618 0 _0466_
rlabel metal1 39054 37230 39054 37230 0 _0467_
rlabel metal1 38778 36890 38778 36890 0 _0468_
rlabel metal1 39606 37366 39606 37366 0 _0469_
rlabel metal1 37720 35530 37720 35530 0 _0470_
rlabel metal1 43470 28458 43470 28458 0 _0471_
rlabel metal2 45218 29172 45218 29172 0 _0472_
rlabel metal1 47840 25942 47840 25942 0 _0473_
rlabel metal1 43286 33490 43286 33490 0 _0474_
rlabel metal2 43010 32878 43010 32878 0 _0475_
rlabel metal1 39238 33898 39238 33898 0 _0476_
rlabel metal1 37398 35020 37398 35020 0 _0477_
rlabel metal1 49358 32436 49358 32436 0 _0478_
rlabel metal1 44574 37910 44574 37910 0 _0479_
rlabel metal1 37628 33898 37628 33898 0 _0480_
rlabel metal1 37582 35088 37582 35088 0 _0481_
rlabel metal1 37628 34034 37628 34034 0 _0482_
rlabel metal1 36892 33422 36892 33422 0 _0483_
rlabel metal1 36984 33286 36984 33286 0 _0484_
rlabel metal1 43470 30702 43470 30702 0 _0485_
rlabel metal1 44804 28186 44804 28186 0 _0486_
rlabel metal2 45402 27642 45402 27642 0 _0487_
rlabel metal2 44850 27132 44850 27132 0 _0488_
rlabel metal1 47518 25874 47518 25874 0 _0489_
rlabel metal1 51290 24718 51290 24718 0 _0490_
rlabel metal1 48484 26962 48484 26962 0 _0491_
rlabel metal1 48806 27574 48806 27574 0 _0492_
rlabel metal1 48024 28050 48024 28050 0 _0493_
rlabel metal2 58098 27812 58098 27812 0 _0494_
rlabel metal1 52946 30600 52946 30600 0 _0495_
rlabel metal2 51934 31892 51934 31892 0 _0496_
rlabel metal2 52578 30396 52578 30396 0 _0497_
rlabel metal2 51014 32062 51014 32062 0 _0498_
rlabel metal1 51934 31858 51934 31858 0 _0499_
rlabel metal1 53130 31858 53130 31858 0 _0500_
rlabel metal2 54510 32708 54510 32708 0 _0501_
rlabel metal2 51750 44166 51750 44166 0 _0502_
rlabel metal1 52808 44234 52808 44234 0 _0503_
rlabel metal1 42412 44234 42412 44234 0 _0504_
rlabel metal1 43976 44982 43976 44982 0 _0505_
rlabel metal1 40112 40902 40112 40902 0 _0506_
rlabel metal2 40802 41990 40802 41990 0 _0507_
rlabel metal2 32982 40188 32982 40188 0 _0508_
rlabel metal2 32338 40494 32338 40494 0 _0509_
rlabel metal2 29302 35836 29302 35836 0 _0510_
rlabel metal2 29854 37842 29854 37842 0 _0511_
rlabel metal2 29118 40868 29118 40868 0 _0512_
rlabel metal1 33212 41106 33212 41106 0 _0513_
rlabel metal2 33718 41922 33718 41922 0 _0514_
rlabel metal1 44620 42194 44620 42194 0 _0515_
rlabel metal2 45770 44642 45770 44642 0 _0516_
rlabel metal2 50554 45050 50554 45050 0 _0517_
rlabel metal2 43378 42364 43378 42364 0 _0518_
rlabel metal1 44160 42330 44160 42330 0 _0519_
rlabel metal2 33534 35700 33534 35700 0 _0520_
rlabel metal2 34086 35836 34086 35836 0 _0521_
rlabel metal1 33856 38930 33856 38930 0 _0522_
rlabel metal1 30544 38318 30544 38318 0 _0523_
rlabel metal1 31004 38522 31004 38522 0 _0524_
rlabel metal2 33534 39678 33534 39678 0 _0525_
rlabel metal1 34592 41514 34592 41514 0 _0526_
rlabel metal1 35604 40698 35604 40698 0 _0527_
rlabel metal1 33626 41004 33626 41004 0 _0528_
rlabel metal1 34454 41242 34454 41242 0 _0529_
rlabel metal1 36018 41684 36018 41684 0 _0530_
rlabel metal2 45586 42500 45586 42500 0 _0531_
rlabel metal1 46782 42568 46782 42568 0 _0532_
rlabel metal2 53038 44642 53038 44642 0 _0533_
rlabel metal1 55384 44370 55384 44370 0 _0534_
rlabel metal1 53176 42330 53176 42330 0 _0535_
rlabel metal1 53728 42874 53728 42874 0 _0536_
rlabel metal2 50370 43962 50370 43962 0 _0537_
rlabel metal1 50830 43962 50830 43962 0 _0538_
rlabel metal2 50922 45220 50922 45220 0 _0539_
rlabel metal2 51566 44336 51566 44336 0 _0540_
rlabel metal1 54326 43962 54326 43962 0 _0541_
rlabel metal1 56304 35054 56304 35054 0 _0542_
rlabel metal1 49036 42670 49036 42670 0 _0543_
rlabel metal1 49910 42874 49910 42874 0 _0544_
rlabel metal1 51175 43214 51175 43214 0 _0545_
rlabel metal1 51612 34510 51612 34510 0 _0546_
rlabel metal2 54510 34170 54510 34170 0 _0547_
rlabel metal2 54234 33796 54234 33796 0 _0548_
rlabel metal2 54050 33796 54050 33796 0 _0549_
rlabel metal2 53774 30022 53774 30022 0 _0550_
rlabel metal1 52762 32912 52762 32912 0 _0551_
rlabel metal2 52946 32708 52946 32708 0 _0552_
rlabel metal2 52394 34068 52394 34068 0 _0553_
rlabel metal1 52532 34442 52532 34442 0 _0554_
rlabel metal1 53314 33388 53314 33388 0 _0555_
rlabel metal2 53406 33932 53406 33932 0 _0556_
rlabel metal2 53130 32581 53130 32581 0 _0557_
rlabel metal2 53590 33762 53590 33762 0 _0558_
rlabel metal2 54050 41820 54050 41820 0 _0559_
rlabel metal1 54924 42874 54924 42874 0 _0560_
rlabel metal1 47656 39406 47656 39406 0 _0561_
rlabel metal1 49266 39542 49266 39542 0 _0562_
rlabel metal2 42366 41786 42366 41786 0 _0563_
rlabel metal1 43424 41582 43424 41582 0 _0564_
rlabel metal1 35512 39066 35512 39066 0 _0565_
rlabel metal2 36110 39814 36110 39814 0 _0566_
rlabel metal2 32246 38522 32246 38522 0 _0567_
rlabel metal1 33212 38318 33212 38318 0 _0568_
rlabel metal2 47058 30957 47058 30957 0 _0569_
rlabel metal1 33534 33626 33534 33626 0 _0570_
rlabel metal1 33120 34170 33120 34170 0 _0571_
rlabel metal1 38364 38930 38364 38930 0 _0572_
rlabel metal1 33948 38862 33948 38862 0 _0573_
rlabel metal2 34086 39780 34086 39780 0 _0574_
rlabel metal2 43930 40460 43930 40460 0 _0575_
rlabel metal1 44804 41650 44804 41650 0 _0576_
rlabel metal1 46322 41684 46322 41684 0 _0577_
rlabel metal2 51290 42432 51290 42432 0 _0578_
rlabel metal1 55062 43180 55062 43180 0 _0579_
rlabel metal2 55338 43486 55338 43486 0 _0580_
rlabel metal1 56488 35122 56488 35122 0 _0581_
rlabel metal2 56258 32708 56258 32708 0 _0582_
rlabel metal1 55568 33082 55568 33082 0 _0583_
rlabel metal1 56028 34510 56028 34510 0 _0584_
rlabel metal2 56074 34170 56074 34170 0 _0585_
rlabel metal2 55982 34442 55982 34442 0 _0586_
rlabel metal1 54096 32538 54096 32538 0 _0587_
rlabel metal1 54556 33082 54556 33082 0 _0588_
rlabel metal2 36938 39100 36938 39100 0 _0589_
rlabel metal1 36800 38726 36800 38726 0 _0590_
rlabel metal1 38640 38386 38640 38386 0 _0591_
rlabel metal1 40020 39406 40020 39406 0 _0592_
rlabel metal2 34454 39168 34454 39168 0 _0593_
rlabel metal1 37300 40018 37300 40018 0 _0594_
rlabel metal2 38134 39644 38134 39644 0 _0595_
rlabel metal2 38870 39746 38870 39746 0 _0596_
rlabel metal2 46690 40188 46690 40188 0 _0597_
rlabel metal1 42642 41072 42642 41072 0 _0598_
rlabel metal1 43838 41004 43838 41004 0 _0599_
rlabel metal1 45310 41038 45310 41038 0 _0600_
rlabel metal1 55154 41072 55154 41072 0 _0601_
rlabel metal1 55936 41242 55936 41242 0 _0602_
rlabel metal1 51152 40902 51152 40902 0 _0603_
rlabel metal1 54464 41718 54464 41718 0 _0604_
rlabel metal1 57178 41650 57178 41650 0 _0605_
rlabel metal1 53774 40698 53774 40698 0 _0606_
rlabel metal2 54786 42534 54786 42534 0 _0607_
rlabel metal1 56810 42806 56810 42806 0 _0608_
rlabel metal1 57270 33626 57270 33626 0 _0609_
rlabel metal1 57408 34374 57408 34374 0 _0610_
rlabel metal1 57687 34714 57687 34714 0 _0611_
rlabel metal1 56672 33966 56672 33966 0 _0612_
rlabel metal1 53222 34000 53222 34000 0 _0613_
rlabel metal2 53038 30702 53038 30702 0 _0614_
rlabel metal2 52026 40698 52026 40698 0 _0615_
rlabel metal1 54188 40630 54188 40630 0 _0616_
rlabel metal1 57040 40018 57040 40018 0 _0617_
rlabel metal1 39560 38182 39560 38182 0 _0618_
rlabel viali 42279 39406 42279 39406 0 _0619_
rlabel metal1 41108 39406 41108 39406 0 _0620_
rlabel metal1 41170 39304 41170 39304 0 _0621_
rlabel metal1 42458 40018 42458 40018 0 _0622_
rlabel metal1 43608 40018 43608 40018 0 _0623_
rlabel metal2 36754 37740 36754 37740 0 _0624_
rlabel metal1 36340 36006 36340 36006 0 _0625_
rlabel metal1 35650 36686 35650 36686 0 _0626_
rlabel metal1 36340 36890 36340 36890 0 _0627_
rlabel metal2 39238 37026 39238 37026 0 _0628_
rlabel metal1 44804 40154 44804 40154 0 _0629_
rlabel metal1 45770 40596 45770 40596 0 _0630_
rlabel metal1 54970 40052 54970 40052 0 _0631_
rlabel metal1 54004 40154 54004 40154 0 _0632_
rlabel metal2 54878 40154 54878 40154 0 _0633_
rlabel metal1 55338 39916 55338 39916 0 _0634_
rlabel metal1 57224 40154 57224 40154 0 _0635_
rlabel metal1 57270 32844 57270 32844 0 _0636_
rlabel metal2 56442 32198 56442 32198 0 _0637_
rlabel metal1 57224 32538 57224 32538 0 _0638_
rlabel metal2 57546 33286 57546 33286 0 _0639_
rlabel metal1 58052 32946 58052 32946 0 _0640_
rlabel metal1 58144 32742 58144 32742 0 _0641_
rlabel metal1 56672 31314 56672 31314 0 _0642_
rlabel metal2 57178 30906 57178 30906 0 _0643_
rlabel metal2 48346 38726 48346 38726 0 _0644_
rlabel metal2 55798 39236 55798 39236 0 _0645_
rlabel metal2 39790 38148 39790 38148 0 _0646_
rlabel metal2 41078 38692 41078 38692 0 _0647_
rlabel metal1 44942 39406 44942 39406 0 _0648_
rlabel metal2 42734 40018 42734 40018 0 _0649_
rlabel metal1 43378 39508 43378 39508 0 _0650_
rlabel metal1 44666 39508 44666 39508 0 _0651_
rlabel metal1 46506 39542 46506 39542 0 _0652_
rlabel metal2 56534 39100 56534 39100 0 _0653_
rlabel metal1 53773 39406 53773 39406 0 _0654_
rlabel metal1 56258 38862 56258 38862 0 _0655_
rlabel metal2 56902 39236 56902 39236 0 _0656_
rlabel metal1 58282 39270 58282 39270 0 _0657_
rlabel metal1 57592 30906 57592 30906 0 _0658_
rlabel metal1 58006 31926 58006 31926 0 _0659_
rlabel metal1 57454 27540 57454 27540 0 _0660_
rlabel metal2 40066 37026 40066 37026 0 _0661_
rlabel metal1 40250 37196 40250 37196 0 _0662_
rlabel metal1 43010 38386 43010 38386 0 _0663_
rlabel metal1 44068 38454 44068 38454 0 _0664_
rlabel metal1 44666 36210 44666 36210 0 _0665_
rlabel metal1 42642 38964 42642 38964 0 _0666_
rlabel metal1 43700 38862 43700 38862 0 _0667_
rlabel metal1 45172 38794 45172 38794 0 _0668_
rlabel metal2 53222 38080 53222 38080 0 _0669_
rlabel metal1 53590 38964 53590 38964 0 _0670_
rlabel metal1 52946 38386 52946 38386 0 _0671_
rlabel metal1 55200 37774 55200 37774 0 _0672_
rlabel metal2 56350 37638 56350 37638 0 _0673_
rlabel metal1 54142 38522 54142 38522 0 _0674_
rlabel metal1 55430 38386 55430 38386 0 _0675_
rlabel metal1 56488 37774 56488 37774 0 _0676_
rlabel metal2 57224 29852 57224 29852 0 _0677_
rlabel metal1 53682 30260 53682 30260 0 _0678_
rlabel metal1 56902 29648 56902 29648 0 _0679_
rlabel metal2 57730 36924 57730 36924 0 _0680_
rlabel metal1 48162 37808 48162 37808 0 _0681_
rlabel metal1 49864 37842 49864 37842 0 _0682_
rlabel metal2 42642 37638 42642 37638 0 _0683_
rlabel metal2 43378 37468 43378 37468 0 _0684_
rlabel metal2 43746 37604 43746 37604 0 _0685_
rlabel metal1 50002 37774 50002 37774 0 _0686_
rlabel metal1 52210 37774 52210 37774 0 _0687_
rlabel metal2 56166 37026 56166 37026 0 _0688_
rlabel metal2 53682 35462 53682 35462 0 _0689_
rlabel metal1 55890 35564 55890 35564 0 _0690_
rlabel metal1 56902 35802 56902 35802 0 _0691_
rlabel metal1 56994 36006 56994 36006 0 _0692_
rlabel metal1 57500 28526 57500 28526 0 _0693_
rlabel metal1 55154 30702 55154 30702 0 _0694_
rlabel metal2 57086 30362 57086 30362 0 _0695_
rlabel metal1 57684 28594 57684 28594 0 _0696_
rlabel metal2 57270 28186 57270 28186 0 _0697_
rlabel metal1 57914 27914 57914 27914 0 _0698_
rlabel metal2 57730 27676 57730 27676 0 _0699_
rlabel metal1 53958 27370 53958 27370 0 _0700_
rlabel metal1 50002 26350 50002 26350 0 _0701_
rlabel metal1 50462 26928 50462 26928 0 _0702_
rlabel metal2 50554 26282 50554 26282 0 _0703_
rlabel metal1 50186 27574 50186 27574 0 _0704_
rlabel metal1 51980 27642 51980 27642 0 _0705_
rlabel metal2 50370 38522 50370 38522 0 _0706_
rlabel metal2 51106 38726 51106 38726 0 _0707_
rlabel metal1 46276 36278 46276 36278 0 _0708_
rlabel metal1 43608 36210 43608 36210 0 _0709_
rlabel metal2 49266 36550 49266 36550 0 _0710_
rlabel metal2 51198 38658 51198 38658 0 _0711_
rlabel metal2 52762 37434 52762 37434 0 _0712_
rlabel metal2 46690 35258 46690 35258 0 _0713_
rlabel metal1 51359 35666 51359 35666 0 _0714_
rlabel metal1 48898 36006 48898 36006 0 _0715_
rlabel metal1 50324 35666 50324 35666 0 _0716_
rlabel metal1 51566 35564 51566 35564 0 _0717_
rlabel metal1 52026 35564 52026 35564 0 _0718_
rlabel metal1 53728 35598 53728 35598 0 _0719_
rlabel metal2 50370 36346 50370 36346 0 _0720_
rlabel metal2 50830 35530 50830 35530 0 _0721_
rlabel metal2 48346 35326 48346 35326 0 _0722_
rlabel metal1 51106 33932 51106 33932 0 _0723_
rlabel metal2 52394 30396 52394 30396 0 _0724_
rlabel metal2 51934 29852 51934 29852 0 _0725_
rlabel metal1 52946 29138 52946 29138 0 _0726_
rlabel metal2 53498 28730 53498 28730 0 _0727_
rlabel metal1 53544 28186 53544 28186 0 _0728_
rlabel metal1 48024 37230 48024 37230 0 _0729_
rlabel metal2 49174 36890 49174 36890 0 _0730_
rlabel metal1 49680 36686 49680 36686 0 _0731_
rlabel via1 53682 36142 53682 36142 0 _0732_
rlabel metal1 54142 37196 54142 37196 0 _0733_
rlabel metal2 54878 36890 54878 36890 0 _0734_
rlabel metal2 55154 36346 55154 36346 0 _0735_
rlabel metal1 55384 36006 55384 36006 0 _0736_
rlabel metal1 52808 36686 52808 36686 0 _0737_
rlabel metal2 52854 36380 52854 36380 0 _0738_
rlabel metal1 53130 36244 53130 36244 0 _0739_
rlabel metal2 54786 28781 54786 28781 0 _0740_
rlabel metal2 55522 29308 55522 29308 0 _0741_
rlabel metal2 54878 28764 54878 28764 0 _0742_
rlabel metal2 54418 28900 54418 28900 0 _0743_
rlabel via1 53695 28526 53695 28526 0 _0744_
rlabel metal2 54142 28220 54142 28220 0 _0745_
rlabel metal2 53958 27914 53958 27914 0 _0746_
rlabel metal1 53728 29614 53728 29614 0 _0747_
rlabel metal2 53314 28186 53314 28186 0 _0748_
rlabel metal2 54326 26996 54326 26996 0 _0749_
rlabel metal2 55062 27166 55062 27166 0 _0750_
rlabel metal2 54694 26758 54694 26758 0 _0751_
rlabel metal2 55982 29580 55982 29580 0 _0752_
rlabel metal2 55614 28458 55614 28458 0 _0753_
rlabel metal2 55890 27642 55890 27642 0 _0754_
rlabel metal2 55154 27166 55154 27166 0 _0755_
rlabel metal1 55338 26928 55338 26928 0 _0756_
rlabel metal2 54786 27200 54786 27200 0 _0757_
rlabel metal1 53084 27302 53084 27302 0 _0758_
rlabel metal2 48254 32640 48254 32640 0 _0759_
rlabel metal1 48484 33082 48484 33082 0 _0760_
rlabel metal2 51106 33184 51106 33184 0 _0761_
rlabel metal1 49220 31178 49220 31178 0 _0762_
rlabel metal1 50968 31450 50968 31450 0 _0763_
rlabel metal1 49956 32334 49956 32334 0 _0764_
rlabel metal2 49818 32708 49818 32708 0 _0765_
rlabel metal1 50232 33082 50232 33082 0 _0766_
rlabel metal2 49818 33252 49818 33252 0 _0767_
rlabel metal2 52210 32198 52210 32198 0 _0768_
rlabel metal1 51474 32538 51474 32538 0 _0769_
rlabel metal1 51934 34000 51934 34000 0 _0770_
rlabel metal2 52026 33694 52026 33694 0 _0771_
rlabel metal2 50278 33660 50278 33660 0 _0772_
rlabel metal1 49772 33286 49772 33286 0 _0773_
rlabel metal2 48162 32096 48162 32096 0 _0774_
rlabel metal2 47610 31178 47610 31178 0 _0775_
rlabel metal1 46506 30736 46506 30736 0 _0776_
rlabel metal1 47196 27574 47196 27574 0 _0777_
rlabel metal2 51658 27489 51658 27489 0 _0778_
rlabel metal2 50646 27744 50646 27744 0 _0779_
rlabel metal1 51290 27642 51290 27642 0 _0780_
rlabel metal2 50370 25670 50370 25670 0 _0781_
rlabel metal2 51198 27404 51198 27404 0 _0782_
rlabel via2 48990 28067 48990 28067 0 _0783_
rlabel metal1 49404 27846 49404 27846 0 _0784_
rlabel metal2 48806 28492 48806 28492 0 _0785_
rlabel metal1 49956 27982 49956 27982 0 _0786_
rlabel metal1 46598 30260 46598 30260 0 _0787_
rlabel metal2 46414 30736 46414 30736 0 _0788_
rlabel metal1 46598 29818 46598 29818 0 _0789_
rlabel metal2 50278 29002 50278 29002 0 _0790_
rlabel metal2 46506 28560 46506 28560 0 _0791_
rlabel metal2 46138 27914 46138 27914 0 _0792_
rlabel metal1 46046 28186 46046 28186 0 _0793_
rlabel metal1 46598 27438 46598 27438 0 _0794_
rlabel metal1 46506 27642 46506 27642 0 _0795_
rlabel metal1 49450 28084 49450 28084 0 _0796_
rlabel metal2 50554 27404 50554 27404 0 _0797_
rlabel metal1 51474 26928 51474 26928 0 _0798_
rlabel metal1 49496 20910 49496 20910 0 clknet_0_net12
rlabel metal1 33396 29546 33396 29546 0 clknet_0_net8
rlabel metal2 47334 21597 47334 21597 0 clknet_1_0__leaf_net12
rlabel metal1 33212 26894 33212 26894 0 clknet_1_0__leaf_net8
rlabel metal1 51198 25330 51198 25330 0 clknet_1_1__leaf_net12
rlabel metal2 34178 30464 34178 30464 0 clknet_1_1__leaf_net8
rlabel metal2 57362 28526 57362 28526 0 count2\[0\]
rlabel metal2 52302 27438 52302 27438 0 count2\[1\]
rlabel metal1 45126 26350 45126 26350 0 count2\[2\]
rlabel metal2 48346 24820 48346 24820 0 count2\[3\]
rlabel metal1 47886 22032 47886 22032 0 count2\[4\]
rlabel metal1 46828 24786 46828 24786 0 count2\[5\]
rlabel metal2 37214 24038 37214 24038 0 count\[0\]
rlabel metal1 38410 27642 38410 27642 0 count\[1\]
rlabel metal1 39146 24072 39146 24072 0 count\[2\]
rlabel metal2 40342 23970 40342 23970 0 count\[3\]
rlabel metal2 37398 22848 37398 22848 0 count\[4\]
rlabel metal1 39560 23698 39560 23698 0 count\[5\]
rlabel metal1 58420 56678 58420 56678 0 net1
rlabel metal1 35742 22066 35742 22066 0 net10
rlabel metal2 43194 30702 43194 30702 0 net11
rlabel metal2 48806 24242 48806 24242 0 net12
rlabel metal2 41078 33728 41078 33728 0 net13
rlabel metal2 39790 24004 39790 24004 0 net14
rlabel metal1 32338 2618 32338 2618 0 net2
rlabel metal1 1886 2618 1886 2618 0 net3
rlabel metal2 1978 57018 1978 57018 0 net4
rlabel metal1 54970 22406 54970 22406 0 net5
rlabel metal1 55338 25398 55338 25398 0 net6
rlabel metal2 2438 28560 2438 28560 0 net7
rlabel metal1 32890 30056 32890 30056 0 net8
rlabel metal2 32982 32096 32982 32096 0 net9
rlabel metal2 1610 1870 1610 1870 0 sel
rlabel metal1 1472 57426 1472 57426 0 user_clock2
rlabel metal2 2070 56406 2070 56406 0 wb_clk_i
rlabel metal1 58466 2346 58466 2346 0 wb_rst_i
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
