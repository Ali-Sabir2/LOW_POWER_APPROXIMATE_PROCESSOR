VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mult_asic_16x16
  CLASS BLOCK ;
  FOREIGN mult_asic_16x16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN A_PAD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 332.640 4.000 333.200 ;
    END
  END A_PAD
  PIN B_PAD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 1.000 333.200 4.000 ;
    END
  END B_PAD
  PIN P0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END P0
  PIN P1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 496.000 165.200 499.000 ;
    END
  END P1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.680 23.840 482.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.680 177.440 482.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.680 331.040 482.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.680 484.640 482.160 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.720 31.530 492.800 33.130 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.720 184.710 492.800 186.310 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.720 337.890 492.800 339.490 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 25.540 15.680 27.140 482.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 179.140 15.680 180.740 482.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 332.740 15.680 334.340 482.160 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 486.340 15.680 487.940 482.160 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.720 34.830 492.800 36.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.720 188.010 492.800 189.610 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 6.720 341.190 492.800 342.790 ;
    END
  END VSS
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 496.000 497.840 499.000 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 164.640 499.000 165.200 ;
    END
  END rst
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 492.800 482.460 ;
      LAYER Metal2 ;
        RECT 0.140 495.700 164.340 496.000 ;
        RECT 165.500 495.700 496.980 496.000 ;
        RECT 0.140 4.300 497.700 495.700 ;
        RECT 0.860 4.000 332.340 4.300 ;
        RECT 333.500 4.000 497.700 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 333.500 497.750 487.620 ;
        RECT 0.090 332.340 0.700 333.500 ;
        RECT 4.300 332.340 497.750 333.500 ;
        RECT 0.090 165.500 497.750 332.340 ;
        RECT 0.090 164.340 495.700 165.500 ;
        RECT 0.090 9.100 497.750 164.340 ;
      LAYER Metal4 ;
        RECT 29.260 25.290 175.540 456.870 ;
        RECT 177.740 25.290 178.840 456.870 ;
        RECT 181.040 25.290 329.140 456.870 ;
        RECT 331.340 25.290 332.440 456.870 ;
        RECT 334.640 25.290 479.220 456.870 ;
      LAYER Metal5 ;
        RECT 29.180 343.290 479.300 343.780 ;
        RECT 29.180 339.990 479.300 340.690 ;
        RECT 29.180 190.110 479.300 337.390 ;
        RECT 29.180 186.810 479.300 187.510 ;
        RECT 29.180 36.930 479.300 184.210 ;
        RECT 29.180 33.630 479.300 34.330 ;
        RECT 29.180 25.260 479.300 31.030 ;
  END
END mult_asic_16x16
END LIBRARY

