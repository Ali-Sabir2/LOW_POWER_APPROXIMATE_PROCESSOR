module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vss,
    vdd,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vss;
 input vdd;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire net73;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net74;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net75;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net146;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net147;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net148;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net149;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net150;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net151;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire \mprj.PS_R1_inst1.LUT_inst1.i0 ;
 wire \mprj.PS_R1_inst1.LUT_inst1.i1 ;
 wire \mprj.PS_R1_inst1.LUT_inst1.i3 ;
 wire \mprj.PS_R1_inst1.LUT_inst1.i4 ;
 wire \mprj.PS_R1_inst1.LUT_inst10.I0 ;
 wire \mprj.PS_R1_inst1.LUT_inst10.I1 ;
 wire \mprj.PS_R1_inst1.LUT_inst11.I1 ;
 wire \mprj.PS_R1_inst1.LUT_inst12.I1 ;
 wire \mprj.PS_R1_inst1.LUT_inst13.I1 ;
 wire \mprj.PS_R1_inst1.LUT_inst14.I1 ;
 wire \mprj.PS_R1_inst1.LUT_inst15.I1 ;
 wire \mprj.PS_R1_inst1.LUT_inst2.I1 ;
 wire \mprj.PS_R1_inst1.LUT_inst3.I1 ;
 wire \mprj.PS_R1_inst1.LUT_inst4.I1 ;
 wire \mprj.PS_R1_inst1.LUT_inst5.I1 ;
 wire \mprj.PS_R1_inst1.LUT_inst6.I1 ;
 wire \mprj.PS_R1_inst1.LUT_inst7.I1 ;
 wire \mprj.PS_R1_inst1.LUT_inst8.I1 ;
 wire \mprj.PS_Rx_inst2.LUT_inst1.i3 ;
 wire \mprj.PS_Rx_inst2.LUT_inst1.i4 ;
 wire \mprj.PS_Rx_inst3.LUT_inst1.i3 ;
 wire \mprj.PS_Rx_inst3.LUT_inst1.i4 ;
 wire \mprj.PS_Rx_inst4.LUT_inst1.i3 ;
 wire \mprj.PS_Rx_inst4.LUT_inst1.i4 ;
 wire \mprj.PS_Rx_inst5.LUT_inst1.i3 ;
 wire \mprj.PS_Rx_inst5.LUT_inst1.i4 ;
 wire \mprj.PS_Rx_inst6.LUT_inst1.i3 ;
 wire \mprj.PS_Rx_inst6.LUT_inst1.i4 ;
 wire \mprj.PS_Rx_inst7.LUT_inst1.i3 ;
 wire \mprj.PS_Rx_inst7.LUT_inst1.i4 ;
 wire \mprj.PS_Rx_inst8.LUT_inst1.i3 ;
 wire \mprj.PS_Rx_inst8.LUT_inst1.i4 ;
 wire \mprj.PS_Rx_inst8.carry_inst.O ;
 wire net210;
 wire net211;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;

 gf180mcu_fd_sc_mcu7t5v0__or4_4 _0674_ (.A1(net10),
    .A2(net9),
    .A3(net12),
    .A4(net11),
    .Z(_0032_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0675_ (.A1(net6),
    .A2(net5),
    .A3(net8),
    .ZN(_0033_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0676_ (.A1(net31),
    .A2(net13),
    .A3(net30),
    .A4(_0033_),
    .ZN(_0034_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0677_ (.A1(_0032_),
    .A2(_0034_),
    .ZN(net35),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _0678_ (.I(\mprj.PS_R1_inst1.LUT_inst1.i0 ),
    .ZN(_0035_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0679_ (.A1(net6),
    .A2(net5),
    .ZN(_0036_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0680_ (.A1(net13),
    .A2(net30),
    .ZN(_0037_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0681_ (.A1(net31),
    .A2(_0037_),
    .ZN(_0038_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0682_ (.A1(net7),
    .A2(_0032_),
    .ZN(_0039_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _0683_ (.A1(_0036_),
    .A2(_0038_),
    .A3(_0039_),
    .Z(_0040_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0684_ (.I(net7),
    .ZN(_0041_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0685_ (.A1(_0041_),
    .A2(_0032_),
    .ZN(_0042_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _0686_ (.A1(_0033_),
    .A2(_0038_),
    .A3(_0042_),
    .ZN(_0043_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _0687_ (.I(_0043_),
    .ZN(_0044_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0688_ (.A1(_0036_),
    .A2(_0039_),
    .B(\mprj.PS_R1_inst1.LUT_inst1.i3 ),
    .ZN(_0045_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0689_ (.A1(_0035_),
    .A2(_0040_),
    .B1(_0044_),
    .B2(_0045_),
    .ZN(net36),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0690_ (.I(\mprj.PS_R1_inst1.LUT_inst1.i4 ),
    .Z(_0046_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _0691_ (.I(\mprj.PS_R1_inst1.LUT_inst1.i3 ),
    .ZN(_0047_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0692_ (.A1(_0035_),
    .A2(\mprj.PS_R1_inst1.LUT_inst1.i1 ),
    .B(_0047_),
    .ZN(_0048_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0693_ (.A1(_0046_),
    .A2(_0048_),
    .ZN(_0049_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0694_ (.A1(net8),
    .A2(_0040_),
    .ZN(_0050_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0695_ (.I(_0050_),
    .Z(_0051_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _0696_ (.I(_0046_),
    .ZN(_0052_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _0697_ (.I(\mprj.PS_R1_inst1.LUT_inst1.i1 ),
    .ZN(_0053_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0698_ (.A1(\mprj.PS_R1_inst1.LUT_inst1.i0 ),
    .A2(_0053_),
    .B(\mprj.PS_R1_inst1.LUT_inst1.i3 ),
    .ZN(_0054_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0699_ (.A1(_0052_),
    .A2(_0054_),
    .ZN(_0055_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0700_ (.A1(_0046_),
    .A2(_0043_),
    .ZN(_0056_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _0701_ (.I(net8),
    .ZN(_0057_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0702_ (.I(_0057_),
    .Z(_0058_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0703_ (.I(\mprj.PS_R1_inst1.LUT_inst1.i1 ),
    .Z(_0059_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _0704_ (.A1(_0036_),
    .A2(_0038_),
    .A3(_0039_),
    .ZN(_0060_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0705_ (.A1(_0058_),
    .A2(_0059_),
    .B(_0060_),
    .ZN(_0061_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _0706_ (.A1(_0049_),
    .A2(_0051_),
    .A3(_0055_),
    .B1(_0056_),
    .B2(_0061_),
    .ZN(net47),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0707_ (.I(\mprj.PS_R1_inst1.LUT_inst2.I1 ),
    .Z(_0062_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0708_ (.I(_0062_),
    .Z(_0063_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0709_ (.I(_0060_),
    .Z(_0064_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0710_ (.I(\mprj.PS_Rx_inst2.LUT_inst1.i3 ),
    .Z(_0065_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _0711_ (.A1(_0063_),
    .A2(_0064_),
    .B1(_0043_),
    .B2(_0065_),
    .C(_0051_),
    .ZN(_0066_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _0712_ (.A1(_0052_),
    .A2(_0048_),
    .A3(_0051_),
    .B(_0066_),
    .ZN(net58),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0713_ (.I(\mprj.PS_Rx_inst2.LUT_inst1.i4 ),
    .Z(_0067_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0714_ (.I(_0043_),
    .Z(_0068_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0715_ (.A1(_0067_),
    .A2(_0068_),
    .ZN(_0069_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0716_ (.I(\mprj.PS_R1_inst1.LUT_inst3.I1 ),
    .Z(_0070_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0717_ (.I(_0070_),
    .Z(_0071_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0718_ (.A1(_0058_),
    .A2(_0071_),
    .B(_0064_),
    .ZN(_0072_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0719_ (.A1(_0046_),
    .A2(_0065_),
    .ZN(_0073_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0720_ (.A1(_0046_),
    .A2(_0065_),
    .Z(_0074_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0721_ (.A1(\mprj.PS_Rx_inst2.LUT_inst1.i4 ),
    .A2(_0073_),
    .A3(_0074_),
    .ZN(_0075_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0722_ (.I(_0075_),
    .Z(_0076_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0723_ (.A1(\mprj.PS_R1_inst1.LUT_inst1.i1 ),
    .A2(_0076_),
    .ZN(_0077_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0724_ (.I(\mprj.PS_R1_inst1.LUT_inst1.i0 ),
    .Z(_0078_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _0725_ (.A1(\mprj.PS_R1_inst1.LUT_inst1.i4 ),
    .A2(_0065_),
    .Z(_0079_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0726_ (.A1(\mprj.PS_R1_inst1.LUT_inst1.i4 ),
    .A2(\mprj.PS_Rx_inst2.LUT_inst1.i3 ),
    .ZN(_0080_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0727_ (.I(_0080_),
    .Z(_0081_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0728_ (.A1(_0078_),
    .A2(_0079_),
    .B(_0081_),
    .ZN(_0082_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0729_ (.A1(_0078_),
    .A2(_0067_),
    .B(_0082_),
    .ZN(_0083_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0730_ (.A1(_0046_),
    .A2(_0054_),
    .B1(_0077_),
    .B2(_0083_),
    .ZN(_0084_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _0731_ (.I(_0084_),
    .ZN(_0085_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0732_ (.A1(_0046_),
    .A2(_0048_),
    .ZN(_0086_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _0733_ (.A1(_0052_),
    .A2(_0065_),
    .B1(_0067_),
    .B2(_0078_),
    .ZN(_0087_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _0734_ (.A1(_0086_),
    .A2(_0077_),
    .A3(_0087_),
    .ZN(_0088_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0735_ (.A1(_0085_),
    .A2(_0088_),
    .ZN(_0089_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0736_ (.A1(_0067_),
    .A2(_0089_),
    .B(_0050_),
    .ZN(_0090_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0737_ (.A1(_0067_),
    .A2(_0089_),
    .B(_0090_),
    .ZN(_0091_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0738_ (.A1(_0069_),
    .A2(_0072_),
    .B(_0091_),
    .ZN(net61),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0739_ (.A1(\mprj.PS_Rx_inst3.LUT_inst1.i3 ),
    .A2(_0044_),
    .ZN(_0092_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0740_ (.I(\mprj.PS_R1_inst1.LUT_inst4.I1 ),
    .Z(_0093_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0741_ (.I(_0093_),
    .Z(_0094_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0742_ (.A1(net8),
    .A2(_0094_),
    .B(_0040_),
    .ZN(_0095_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0743_ (.A1(_0065_),
    .A2(_0067_),
    .B(_0059_),
    .ZN(_0096_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0744_ (.A1(_0067_),
    .A2(_0073_),
    .B(_0074_),
    .ZN(_0097_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0745_ (.A1(_0046_),
    .A2(_0065_),
    .B(\mprj.PS_Rx_inst2.LUT_inst1.i4 ),
    .ZN(_0098_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0746_ (.I(_0098_),
    .Z(_0099_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _0747_ (.A1(_0096_),
    .A2(_0097_),
    .B1(_0099_),
    .B2(_0063_),
    .ZN(_0100_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0748_ (.A1(_0063_),
    .A2(_0076_),
    .B(_0100_),
    .ZN(_0101_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0749_ (.A1(_0057_),
    .A2(_0060_),
    .ZN(_0102_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _0750_ (.I(_0102_),
    .Z(_0103_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0751_ (.A1(_0092_),
    .A2(_0095_),
    .B1(_0101_),
    .B2(_0103_),
    .ZN(net62),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0752_ (.I(\mprj.PS_Rx_inst3.LUT_inst1.i4 ),
    .Z(_0104_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0753_ (.A1(_0104_),
    .A2(_0068_),
    .ZN(_0105_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0754_ (.I(\mprj.PS_R1_inst1.LUT_inst5.I1 ),
    .Z(_0106_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0755_ (.I(_0106_),
    .Z(_0107_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0756_ (.A1(_0058_),
    .A2(_0107_),
    .B(_0064_),
    .ZN(_0108_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0757_ (.A1(_0065_),
    .A2(_0067_),
    .B(_0062_),
    .ZN(_0109_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _0758_ (.A1(_0071_),
    .A2(_0099_),
    .B1(_0109_),
    .B2(_0097_),
    .ZN(_0110_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0759_ (.A1(_0071_),
    .A2(_0076_),
    .B(_0110_),
    .ZN(_0111_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _0760_ (.I(_0104_),
    .ZN(_0112_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0761_ (.A1(\mprj.PS_Rx_inst2.LUT_inst1.i4 ),
    .A2(\mprj.PS_Rx_inst3.LUT_inst1.i3 ),
    .ZN(_0113_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _0762_ (.A1(\mprj.PS_Rx_inst2.LUT_inst1.i4 ),
    .A2(\mprj.PS_Rx_inst3.LUT_inst1.i3 ),
    .Z(_0114_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _0763_ (.A1(_0112_),
    .A2(_0113_),
    .A3(_0114_),
    .Z(_0115_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0764_ (.I(_0115_),
    .Z(_0116_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0765_ (.A1(\mprj.PS_Rx_inst3.LUT_inst1.i3 ),
    .A2(_0104_),
    .Z(_0117_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0766_ (.A1(_0078_),
    .A2(_0104_),
    .ZN(_0118_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0767_ (.I(_0113_),
    .Z(_0119_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _0768_ (.A1(_0078_),
    .A2(_0067_),
    .A3(_0117_),
    .B1(_0118_),
    .B2(_0119_),
    .ZN(_0120_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0769_ (.A1(_0059_),
    .A2(_0116_),
    .B(_0120_),
    .ZN(_0121_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0770_ (.A1(_0104_),
    .A2(_0121_),
    .Z(_0122_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0771_ (.A1(_0111_),
    .A2(_0122_),
    .B(_0050_),
    .ZN(_0123_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0772_ (.A1(_0111_),
    .A2(_0122_),
    .B(_0123_),
    .ZN(_0124_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0773_ (.A1(_0105_),
    .A2(_0108_),
    .B(_0124_),
    .ZN(net63),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0774_ (.A1(\mprj.PS_Rx_inst4.LUT_inst1.i3 ),
    .A2(_0068_),
    .ZN(_0125_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0775_ (.I(\mprj.PS_R1_inst1.LUT_inst6.I1 ),
    .Z(_0126_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0776_ (.I(_0126_),
    .Z(_0127_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0777_ (.A1(_0058_),
    .A2(_0127_),
    .B(_0064_),
    .ZN(_0128_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0778_ (.A1(\mprj.PS_Rx_inst2.LUT_inst1.i4 ),
    .A2(\mprj.PS_Rx_inst3.LUT_inst1.i3 ),
    .B(_0104_),
    .ZN(_0129_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0779_ (.I(_0129_),
    .Z(_0130_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0780_ (.A1(_0112_),
    .A2(_0114_),
    .B(_0113_),
    .ZN(_0131_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0781_ (.I(_0131_),
    .Z(_0132_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0782_ (.A1(_0059_),
    .A2(_0117_),
    .B(_0132_),
    .ZN(_0133_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0783_ (.A1(_0063_),
    .A2(_0116_),
    .ZN(_0134_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _0784_ (.A1(_0063_),
    .A2(_0130_),
    .B(_0133_),
    .C(_0134_),
    .ZN(_0135_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _0785_ (.I(\mprj.PS_Rx_inst2.LUT_inst1.i4 ),
    .ZN(_0136_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0786_ (.A1(_0136_),
    .A2(_0079_),
    .B(_0080_),
    .ZN(_0137_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0787_ (.I(_0137_),
    .Z(_0138_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0788_ (.A1(_0094_),
    .A2(_0081_),
    .B(_0099_),
    .ZN(_0139_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0789_ (.A1(_0094_),
    .A2(_0076_),
    .B1(_0138_),
    .B2(_0070_),
    .C(_0139_),
    .ZN(_0140_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0790_ (.A1(_0111_),
    .A2(_0140_),
    .Z(_0141_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0791_ (.A1(_0135_),
    .A2(_0141_),
    .Z(_0142_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0792_ (.A1(_0135_),
    .A2(_0141_),
    .B(_0103_),
    .ZN(_0143_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _0793_ (.A1(_0125_),
    .A2(_0128_),
    .B1(_0142_),
    .B2(_0143_),
    .ZN(net64),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0794_ (.I(\mprj.PS_Rx_inst4.LUT_inst1.i4 ),
    .Z(_0144_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0795_ (.A1(_0144_),
    .A2(_0068_),
    .ZN(_0145_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0796_ (.I(\mprj.PS_R1_inst1.LUT_inst7.I1 ),
    .Z(_0146_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0797_ (.I(_0146_),
    .Z(_0147_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0798_ (.A1(_0058_),
    .A2(_0147_),
    .B(_0064_),
    .ZN(_0148_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0799_ (.A1(\mprj.PS_Rx_inst4.LUT_inst1.i3 ),
    .A2(_0144_),
    .Z(_0149_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0800_ (.A1(_0078_),
    .A2(_0144_),
    .ZN(_0150_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0801_ (.A1(_0104_),
    .A2(\mprj.PS_Rx_inst4.LUT_inst1.i3 ),
    .ZN(_0151_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0802_ (.I(_0151_),
    .Z(_0152_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _0803_ (.A1(_0078_),
    .A2(_0104_),
    .A3(_0149_),
    .B1(_0150_),
    .B2(_0152_),
    .ZN(_0153_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _0804_ (.I(\mprj.PS_Rx_inst4.LUT_inst1.i4 ),
    .ZN(_0154_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _0805_ (.A1(_0104_),
    .A2(\mprj.PS_Rx_inst4.LUT_inst1.i3 ),
    .Z(_0155_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _0806_ (.A1(_0154_),
    .A2(_0151_),
    .A3(_0155_),
    .Z(_0156_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0807_ (.I(_0156_),
    .Z(_0157_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _0808_ (.A1(_0059_),
    .A2(_0157_),
    .B(_0153_),
    .C(_0144_),
    .ZN(_0158_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0809_ (.A1(_0144_),
    .A2(_0153_),
    .B(_0158_),
    .ZN(_0159_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0810_ (.A1(_0070_),
    .A2(_0116_),
    .ZN(_0160_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0811_ (.A1(\mprj.PS_R1_inst1.LUT_inst2.I1 ),
    .A2(_0117_),
    .B(_0132_),
    .ZN(_0161_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _0812_ (.A1(_0070_),
    .A2(_0130_),
    .B(_0160_),
    .C(_0161_),
    .ZN(_0162_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0813_ (.A1(_0106_),
    .A2(_0081_),
    .B(_0099_),
    .ZN(_0163_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0814_ (.A1(_0107_),
    .A2(_0076_),
    .B1(_0138_),
    .B2(_0093_),
    .C(_0163_),
    .ZN(_0164_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _0815_ (.A1(_0140_),
    .A2(_0162_),
    .A3(_0164_),
    .Z(_0165_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0816_ (.A1(_0159_),
    .A2(_0165_),
    .B(_0050_),
    .ZN(_0166_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0817_ (.A1(_0159_),
    .A2(_0165_),
    .B(_0166_),
    .ZN(_0167_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0818_ (.A1(_0145_),
    .A2(_0148_),
    .B(_0167_),
    .ZN(net65),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0819_ (.A1(\mprj.PS_Rx_inst5.LUT_inst1.i3 ),
    .A2(_0044_),
    .ZN(_0168_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0820_ (.I(\mprj.PS_R1_inst1.LUT_inst8.I1 ),
    .Z(_0169_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0821_ (.I(_0169_),
    .Z(_0170_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0822_ (.A1(net8),
    .A2(_0170_),
    .B(_0040_),
    .ZN(_0171_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0823_ (.A1(\mprj.PS_Rx_inst4.LUT_inst1.i4 ),
    .A2(_0155_),
    .ZN(_0172_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0824_ (.I(_0172_),
    .Z(_0173_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0825_ (.A1(_0154_),
    .A2(_0155_),
    .B(_0151_),
    .ZN(_0174_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0826_ (.I(_0174_),
    .Z(_0175_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0827_ (.A1(_0059_),
    .A2(_0149_),
    .B(_0175_),
    .ZN(_0176_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0828_ (.A1(_0062_),
    .A2(_0157_),
    .ZN(_0177_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _0829_ (.A1(_0063_),
    .A2(_0173_),
    .B(_0176_),
    .C(_0177_),
    .ZN(_0178_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0830_ (.A1(_0126_),
    .A2(_0081_),
    .B(_0099_),
    .ZN(_0179_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0831_ (.A1(_0126_),
    .A2(_0076_),
    .B1(_0138_),
    .B2(_0106_),
    .C(_0179_),
    .ZN(_0180_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0832_ (.A1(_0093_),
    .A2(_0119_),
    .B(_0130_),
    .ZN(_0181_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0833_ (.A1(_0093_),
    .A2(_0116_),
    .B1(_0132_),
    .B2(\mprj.PS_R1_inst1.LUT_inst3.I1 ),
    .C(_0181_),
    .ZN(_0182_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _0834_ (.A1(_0164_),
    .A2(_0180_),
    .A3(_0182_),
    .Z(_0183_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0835_ (.A1(_0165_),
    .A2(_0183_),
    .Z(_0184_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0836_ (.A1(_0178_),
    .A2(_0184_),
    .B(_0102_),
    .ZN(_0185_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0837_ (.A1(_0178_),
    .A2(_0184_),
    .B(_0185_),
    .ZN(_0186_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0838_ (.A1(_0168_),
    .A2(_0171_),
    .B(_0186_),
    .ZN(net66),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0839_ (.I(\mprj.PS_Rx_inst5.LUT_inst1.i4 ),
    .Z(_0187_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0840_ (.A1(_0187_),
    .A2(_0068_),
    .ZN(_0188_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0841_ (.I(\mprj.PS_R1_inst1.LUT_inst10.I0 ),
    .Z(_0189_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0842_ (.I(_0189_),
    .Z(_0190_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0843_ (.A1(_0058_),
    .A2(_0190_),
    .B(_0064_),
    .ZN(_0191_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0844_ (.A1(_0070_),
    .A2(_0157_),
    .ZN(_0192_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0845_ (.A1(\mprj.PS_R1_inst1.LUT_inst2.I1 ),
    .A2(_0149_),
    .B(_0175_),
    .ZN(_0193_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _0846_ (.A1(_0071_),
    .A2(_0173_),
    .B(_0192_),
    .C(_0193_),
    .ZN(_0194_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0847_ (.A1(_0146_),
    .A2(_0081_),
    .B(_0099_),
    .ZN(_0195_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0848_ (.A1(_0146_),
    .A2(_0076_),
    .B1(_0138_),
    .B2(_0126_),
    .C(_0195_),
    .ZN(_0196_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0849_ (.A1(_0106_),
    .A2(_0119_),
    .B(_0130_),
    .ZN(_0197_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0850_ (.A1(_0106_),
    .A2(_0116_),
    .B1(_0132_),
    .B2(\mprj.PS_R1_inst1.LUT_inst4.I1 ),
    .C(_0197_),
    .ZN(_0198_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _0851_ (.A1(_0180_),
    .A2(_0196_),
    .A3(_0198_),
    .Z(_0199_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _0852_ (.A1(_0183_),
    .A2(_0194_),
    .A3(_0199_),
    .Z(_0200_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _0853_ (.I(_0187_),
    .ZN(_0201_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _0854_ (.A1(\mprj.PS_Rx_inst4.LUT_inst1.i4 ),
    .A2(\mprj.PS_Rx_inst5.LUT_inst1.i3 ),
    .Z(_0202_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0855_ (.A1(_0201_),
    .A2(_0202_),
    .ZN(_0203_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0856_ (.A1(_0144_),
    .A2(\mprj.PS_Rx_inst5.LUT_inst1.i3 ),
    .B(_0203_),
    .ZN(_0204_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0857_ (.I(_0204_),
    .Z(_0205_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0858_ (.A1(\mprj.PS_Rx_inst5.LUT_inst1.i3 ),
    .A2(_0187_),
    .Z(_0206_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0859_ (.A1(\mprj.PS_R1_inst1.LUT_inst1.i0 ),
    .A2(_0187_),
    .ZN(_0207_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0860_ (.A1(_0144_),
    .A2(\mprj.PS_Rx_inst5.LUT_inst1.i3 ),
    .ZN(_0208_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0861_ (.I(_0208_),
    .Z(_0209_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _0862_ (.A1(_0078_),
    .A2(_0144_),
    .A3(_0206_),
    .B1(_0207_),
    .B2(_0209_),
    .ZN(_0210_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0863_ (.A1(_0059_),
    .A2(_0205_),
    .B(_0210_),
    .ZN(_0211_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0864_ (.A1(_0201_),
    .A2(_0211_),
    .Z(_0212_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0865_ (.A1(_0200_),
    .A2(_0212_),
    .B(_0050_),
    .ZN(_0213_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0866_ (.A1(_0200_),
    .A2(_0212_),
    .B(_0213_),
    .ZN(_0214_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0867_ (.A1(_0188_),
    .A2(_0191_),
    .B(_0214_),
    .ZN(net67),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0868_ (.A1(\mprj.PS_Rx_inst6.LUT_inst1.i3 ),
    .A2(_0068_),
    .ZN(_0215_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0869_ (.I(\mprj.PS_R1_inst1.LUT_inst10.I1 ),
    .Z(_0216_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0870_ (.I(_0216_),
    .Z(_0217_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0871_ (.A1(_0058_),
    .A2(_0217_),
    .B(_0064_),
    .ZN(_0218_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0872_ (.A1(_0187_),
    .A2(_0202_),
    .ZN(_0219_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0873_ (.I(_0219_),
    .Z(_0220_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0874_ (.A1(_0201_),
    .A2(_0202_),
    .B(_0208_),
    .ZN(_0221_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0875_ (.I(_0221_),
    .Z(_0222_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0876_ (.A1(_0059_),
    .A2(_0206_),
    .B(_0222_),
    .ZN(_0223_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0877_ (.A1(_0063_),
    .A2(_0205_),
    .ZN(_0224_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _0878_ (.A1(_0063_),
    .A2(_0220_),
    .B(_0223_),
    .C(_0224_),
    .ZN(_0225_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0879_ (.A1(_0126_),
    .A2(_0119_),
    .B(_0130_),
    .ZN(_0226_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0880_ (.A1(_0126_),
    .A2(_0116_),
    .B1(_0132_),
    .B2(\mprj.PS_R1_inst1.LUT_inst5.I1 ),
    .C(_0226_),
    .ZN(_0227_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0881_ (.A1(\mprj.PS_R1_inst1.LUT_inst8.I1 ),
    .A2(_0080_),
    .B(_0098_),
    .ZN(_0228_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0882_ (.A1(_0169_),
    .A2(_0075_),
    .B1(_0137_),
    .B2(\mprj.PS_R1_inst1.LUT_inst7.I1 ),
    .C(_0228_),
    .ZN(_0229_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _0883_ (.A1(_0196_),
    .A2(_0227_),
    .A3(_0229_),
    .ZN(_0230_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0884_ (.A1(_0093_),
    .A2(_0152_),
    .B(_0173_),
    .ZN(_0231_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0885_ (.A1(_0093_),
    .A2(_0157_),
    .B1(_0175_),
    .B2(\mprj.PS_R1_inst1.LUT_inst3.I1 ),
    .C(_0231_),
    .ZN(_0232_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _0886_ (.A1(_0199_),
    .A2(_0230_),
    .A3(_0232_),
    .Z(_0233_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0887_ (.A1(_0200_),
    .A2(_0233_),
    .Z(_0234_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0888_ (.A1(_0225_),
    .A2(_0234_),
    .Z(_0235_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0889_ (.A1(_0225_),
    .A2(_0234_),
    .B(_0103_),
    .ZN(_0236_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _0890_ (.A1(_0215_),
    .A2(_0218_),
    .B1(_0235_),
    .B2(_0236_),
    .ZN(net37),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0891_ (.I(\mprj.PS_Rx_inst6.LUT_inst1.i4 ),
    .Z(_0237_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0892_ (.A1(_0237_),
    .A2(_0068_),
    .ZN(_0238_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0893_ (.I(\mprj.PS_R1_inst1.LUT_inst11.I1 ),
    .Z(_0239_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0894_ (.I(_0239_),
    .Z(_0240_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0895_ (.A1(_0058_),
    .A2(_0240_),
    .B(_0064_),
    .ZN(_0241_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _0896_ (.I(\mprj.PS_Rx_inst6.LUT_inst1.i4 ),
    .ZN(_0242_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0897_ (.A1(\mprj.PS_Rx_inst6.LUT_inst1.i3 ),
    .A2(_0237_),
    .ZN(_0243_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0898_ (.A1(_0187_),
    .A2(\mprj.PS_Rx_inst6.LUT_inst1.i3 ),
    .ZN(_0244_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0899_ (.A1(_0187_),
    .A2(\mprj.PS_Rx_inst6.LUT_inst1.i3 ),
    .ZN(_0245_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0900_ (.A1(_0242_),
    .A2(_0245_),
    .ZN(_0246_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0901_ (.A1(_0244_),
    .A2(_0246_),
    .ZN(_0247_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0902_ (.I(_0247_),
    .Z(_0248_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _0903_ (.I(_0245_),
    .Z(_0249_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0904_ (.A1(_0078_),
    .A2(_0237_),
    .ZN(_0250_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0905_ (.A1(_0249_),
    .A2(_0250_),
    .ZN(_0251_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0906_ (.A1(_0207_),
    .A2(_0243_),
    .B1(_0248_),
    .B2(_0059_),
    .C(_0251_),
    .ZN(_0252_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0907_ (.A1(_0242_),
    .A2(_0252_),
    .Z(_0253_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0908_ (.A1(_0106_),
    .A2(_0152_),
    .B(_0173_),
    .ZN(_0254_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _0909_ (.A1(_0106_),
    .A2(_0157_),
    .B1(_0175_),
    .B2(\mprj.PS_R1_inst1.LUT_inst4.I1 ),
    .C(_0254_),
    .ZN(_0255_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0910_ (.A1(\mprj.PS_R1_inst1.LUT_inst7.I1 ),
    .A2(_0113_),
    .B(_0129_),
    .ZN(_0256_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0911_ (.A1(\mprj.PS_R1_inst1.LUT_inst7.I1 ),
    .A2(_0115_),
    .B1(_0131_),
    .B2(\mprj.PS_R1_inst1.LUT_inst6.I1 ),
    .C(_0256_),
    .ZN(_0257_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0912_ (.A1(\mprj.PS_R1_inst1.LUT_inst10.I0 ),
    .A2(_0080_),
    .B(_0098_),
    .ZN(_0258_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0913_ (.A1(\mprj.PS_R1_inst1.LUT_inst10.I0 ),
    .A2(_0075_),
    .B1(_0137_),
    .B2(\mprj.PS_R1_inst1.LUT_inst8.I1 ),
    .C(_0258_),
    .ZN(_0259_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _0914_ (.A1(_0229_),
    .A2(_0257_),
    .A3(_0259_),
    .Z(_0260_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _0915_ (.A1(_0230_),
    .A2(_0255_),
    .A3(_0260_),
    .Z(_0261_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0916_ (.A1(_0071_),
    .A2(_0205_),
    .ZN(_0262_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0917_ (.A1(_0062_),
    .A2(_0206_),
    .B(_0222_),
    .ZN(_0263_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _0918_ (.A1(_0071_),
    .A2(_0220_),
    .B(_0262_),
    .C(_0263_),
    .ZN(_0264_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _0919_ (.A1(_0233_),
    .A2(_0261_),
    .A3(_0264_),
    .Z(_0265_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0920_ (.A1(_0253_),
    .A2(_0265_),
    .Z(_0266_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0921_ (.A1(_0253_),
    .A2(_0265_),
    .B(_0103_),
    .ZN(_0267_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _0922_ (.A1(_0238_),
    .A2(_0241_),
    .B1(_0266_),
    .B2(_0267_),
    .ZN(net38),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0923_ (.A1(\mprj.PS_Rx_inst7.LUT_inst1.i3 ),
    .A2(_0068_),
    .ZN(_0268_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0924_ (.I(\mprj.PS_R1_inst1.LUT_inst12.I1 ),
    .Z(_0269_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0925_ (.I(_0269_),
    .Z(_0270_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0926_ (.A1(_0058_),
    .A2(_0270_),
    .B(_0064_),
    .ZN(_0271_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0927_ (.A1(_0093_),
    .A2(_0209_),
    .B(_0220_),
    .ZN(_0272_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0928_ (.A1(_0093_),
    .A2(_0205_),
    .B1(_0222_),
    .B2(\mprj.PS_R1_inst1.LUT_inst3.I1 ),
    .C(_0272_),
    .ZN(_0273_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0929_ (.A1(\mprj.PS_R1_inst1.LUT_inst6.I1 ),
    .A2(_0152_),
    .B(_0172_),
    .ZN(_0274_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0930_ (.A1(\mprj.PS_R1_inst1.LUT_inst6.I1 ),
    .A2(_0156_),
    .B1(_0174_),
    .B2(\mprj.PS_R1_inst1.LUT_inst5.I1 ),
    .C(_0274_),
    .ZN(_0275_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0931_ (.A1(\mprj.PS_R1_inst1.LUT_inst8.I1 ),
    .A2(_0113_),
    .B(_0129_),
    .ZN(_0276_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0932_ (.A1(\mprj.PS_R1_inst1.LUT_inst8.I1 ),
    .A2(_0115_),
    .B1(_0131_),
    .B2(\mprj.PS_R1_inst1.LUT_inst7.I1 ),
    .C(_0276_),
    .ZN(_0277_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0933_ (.A1(\mprj.PS_R1_inst1.LUT_inst10.I1 ),
    .A2(_0081_),
    .B(_0099_),
    .ZN(_0278_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0934_ (.A1(\mprj.PS_R1_inst1.LUT_inst10.I1 ),
    .A2(_0075_),
    .B1(_0138_),
    .B2(\mprj.PS_R1_inst1.LUT_inst10.I0 ),
    .C(_0278_),
    .ZN(_0279_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _0935_ (.A1(_0259_),
    .A2(_0277_),
    .A3(_0279_),
    .Z(_0280_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _0936_ (.A1(_0260_),
    .A2(_0275_),
    .A3(_0280_),
    .ZN(_0281_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _0937_ (.A1(_0261_),
    .A2(_0273_),
    .A3(_0281_),
    .Z(_0282_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0938_ (.A1(\mprj.PS_Rx_inst6.LUT_inst1.i3 ),
    .A2(_0237_),
    .B(\mprj.PS_R1_inst1.LUT_inst1.i1 ),
    .ZN(_0283_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _0939_ (.I(_0283_),
    .ZN(_0284_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0940_ (.A1(\mprj.PS_Rx_inst6.LUT_inst1.i4 ),
    .A2(_0244_),
    .ZN(_0285_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0941_ (.A1(_0245_),
    .A2(_0285_),
    .ZN(_0286_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0942_ (.I(_0286_),
    .Z(_0287_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0943_ (.A1(_0187_),
    .A2(\mprj.PS_Rx_inst6.LUT_inst1.i3 ),
    .B(\mprj.PS_Rx_inst6.LUT_inst1.i4 ),
    .ZN(_0288_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _0944_ (.I(_0288_),
    .Z(_0289_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0945_ (.A1(_0062_),
    .A2(_0289_),
    .ZN(_0290_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0946_ (.A1(_0062_),
    .A2(_0248_),
    .B1(_0284_),
    .B2(_0287_),
    .C(_0290_),
    .ZN(_0291_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _0947_ (.A1(_0265_),
    .A2(_0291_),
    .Z(_0292_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0948_ (.A1(_0282_),
    .A2(_0292_),
    .B(_0050_),
    .ZN(_0293_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0949_ (.A1(_0282_),
    .A2(_0292_),
    .B(_0293_),
    .ZN(_0294_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0950_ (.A1(_0268_),
    .A2(_0271_),
    .B(_0294_),
    .ZN(net39),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0951_ (.I(\mprj.PS_Rx_inst7.LUT_inst1.i4 ),
    .Z(_0295_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0952_ (.A1(_0295_),
    .A2(_0068_),
    .ZN(_0296_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0953_ (.I(\mprj.PS_R1_inst1.LUT_inst13.I1 ),
    .Z(_0297_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0954_ (.I(_0297_),
    .Z(_0298_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0955_ (.A1(_0058_),
    .A2(_0298_),
    .B(_0060_),
    .ZN(_0299_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0956_ (.A1(\mprj.PS_Rx_inst6.LUT_inst1.i3 ),
    .A2(_0237_),
    .B(\mprj.PS_R1_inst1.LUT_inst2.I1 ),
    .ZN(_0300_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0957_ (.I(_0300_),
    .ZN(_0301_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0958_ (.A1(_0070_),
    .A2(_0248_),
    .B1(_0287_),
    .B2(_0301_),
    .ZN(_0302_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0959_ (.A1(_0070_),
    .A2(_0289_),
    .B(_0302_),
    .ZN(_0303_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0960_ (.A1(\mprj.PS_R1_inst1.LUT_inst5.I1 ),
    .A2(_0209_),
    .B(_0219_),
    .ZN(_0304_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0961_ (.A1(_0106_),
    .A2(_0204_),
    .B1(_0221_),
    .B2(\mprj.PS_R1_inst1.LUT_inst4.I1 ),
    .C(_0304_),
    .ZN(_0305_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0962_ (.A1(_0146_),
    .A2(_0151_),
    .B(_0172_),
    .ZN(_0306_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0963_ (.A1(_0146_),
    .A2(_0156_),
    .B1(_0174_),
    .B2(\mprj.PS_R1_inst1.LUT_inst6.I1 ),
    .C(_0306_),
    .ZN(_0307_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0964_ (.A1(\mprj.PS_R1_inst1.LUT_inst10.I0 ),
    .A2(_0119_),
    .B(_0129_),
    .ZN(_0308_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0965_ (.A1(_0189_),
    .A2(_0115_),
    .B1(_0131_),
    .B2(_0169_),
    .C(_0308_),
    .ZN(_0309_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0966_ (.A1(\mprj.PS_R1_inst1.LUT_inst11.I1 ),
    .A2(_0081_),
    .B(_0099_),
    .ZN(_0310_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0967_ (.A1(\mprj.PS_R1_inst1.LUT_inst11.I1 ),
    .A2(_0076_),
    .B1(_0138_),
    .B2(\mprj.PS_R1_inst1.LUT_inst10.I1 ),
    .C(_0310_),
    .ZN(_0311_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_4 _0968_ (.A1(_0279_),
    .A2(_0309_),
    .A3(_0311_),
    .ZN(_0312_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _0969_ (.A1(_0280_),
    .A2(_0307_),
    .A3(_0312_),
    .Z(_0313_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _0970_ (.A1(_0281_),
    .A2(_0305_),
    .A3(_0313_),
    .ZN(_0314_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _0971_ (.A1(_0282_),
    .A2(_0303_),
    .A3(_0314_),
    .Z(_0315_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0972_ (.A1(_0237_),
    .A2(\mprj.PS_Rx_inst7.LUT_inst1.i3 ),
    .ZN(_0316_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0973_ (.A1(_0237_),
    .A2(\mprj.PS_Rx_inst7.LUT_inst1.i3 ),
    .ZN(_0317_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0974_ (.A1(_0295_),
    .A2(_0317_),
    .ZN(_0318_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0975_ (.A1(_0316_),
    .A2(_0318_),
    .Z(_0319_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0976_ (.I(_0319_),
    .Z(_0320_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0977_ (.A1(\mprj.PS_Rx_inst7.LUT_inst1.i3 ),
    .A2(_0295_),
    .ZN(_0321_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _0978_ (.I(_0295_),
    .ZN(_0322_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0979_ (.I(_0316_),
    .Z(_0323_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0980_ (.A1(_0035_),
    .A2(_0322_),
    .B(_0323_),
    .ZN(_0324_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0981_ (.A1(_0059_),
    .A2(_0320_),
    .B1(_0321_),
    .B2(_0250_),
    .C(_0324_),
    .ZN(_0325_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _0982_ (.A1(_0295_),
    .A2(_0325_),
    .Z(_0326_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0983_ (.A1(_0315_),
    .A2(_0326_),
    .Z(_0327_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0984_ (.A1(_0315_),
    .A2(_0326_),
    .B(_0102_),
    .ZN(_0328_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _0985_ (.A1(_0296_),
    .A2(_0299_),
    .B1(_0327_),
    .B2(_0328_),
    .ZN(net40),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0986_ (.A1(\mprj.PS_Rx_inst8.LUT_inst1.i3 ),
    .A2(_0044_),
    .ZN(_0329_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0987_ (.I(\mprj.PS_R1_inst1.LUT_inst14.I1 ),
    .Z(_0330_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0988_ (.I(_0330_),
    .Z(_0331_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0989_ (.A1(net8),
    .A2(_0331_),
    .B(_0040_),
    .ZN(_0332_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0990_ (.A1(_0237_),
    .A2(\mprj.PS_Rx_inst7.LUT_inst1.i3 ),
    .B(_0295_),
    .ZN(_0333_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _0991_ (.I(_0333_),
    .Z(_0334_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0992_ (.A1(_0295_),
    .A2(_0317_),
    .ZN(_0335_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0993_ (.A1(_0316_),
    .A2(_0335_),
    .ZN(_0336_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _0994_ (.I(_0336_),
    .Z(_0337_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0995_ (.A1(_0053_),
    .A2(_0321_),
    .ZN(_0338_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0996_ (.A1(_0062_),
    .A2(_0320_),
    .B1(_0337_),
    .B2(_0338_),
    .ZN(_0339_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0997_ (.A1(_0063_),
    .A2(_0334_),
    .B(_0339_),
    .ZN(_0340_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0998_ (.A1(\mprj.PS_R1_inst1.LUT_inst4.I1 ),
    .A2(_0245_),
    .B(_0288_),
    .ZN(_0341_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0999_ (.A1(_0093_),
    .A2(_0247_),
    .B1(_0286_),
    .B2(\mprj.PS_R1_inst1.LUT_inst3.I1 ),
    .C(_0341_),
    .ZN(_0342_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1000_ (.A1(_0126_),
    .A2(_0208_),
    .B(_0219_),
    .ZN(_0343_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1001_ (.A1(_0126_),
    .A2(_0204_),
    .B1(_0221_),
    .B2(\mprj.PS_R1_inst1.LUT_inst5.I1 ),
    .C(_0343_),
    .ZN(_0344_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1002_ (.A1(_0169_),
    .A2(_0152_),
    .B(_0173_),
    .ZN(_0345_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1003_ (.A1(_0169_),
    .A2(_0156_),
    .B1(_0175_),
    .B2(_0146_),
    .C(_0345_),
    .ZN(_0346_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1004_ (.A1(\mprj.PS_R1_inst1.LUT_inst10.I1 ),
    .A2(_0119_),
    .B(_0129_),
    .ZN(_0347_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1005_ (.A1(_0216_),
    .A2(_0115_),
    .B1(_0131_),
    .B2(_0189_),
    .C(_0347_),
    .ZN(_0348_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1006_ (.A1(\mprj.PS_R1_inst1.LUT_inst12.I1 ),
    .A2(_0081_),
    .B(_0099_),
    .ZN(_0349_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1007_ (.A1(_0269_),
    .A2(_0076_),
    .B1(_0138_),
    .B2(_0239_),
    .C(_0349_),
    .ZN(_0350_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1008_ (.A1(_0311_),
    .A2(_0348_),
    .A3(_0350_),
    .Z(_0351_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1009_ (.A1(_0312_),
    .A2(_0346_),
    .A3(_0351_),
    .Z(_0352_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1010_ (.A1(_0313_),
    .A2(_0344_),
    .A3(_0352_),
    .ZN(_0353_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1011_ (.A1(_0314_),
    .A2(_0342_),
    .A3(_0353_),
    .Z(_0354_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _1012_ (.A1(_0315_),
    .A2(_0354_),
    .ZN(_0355_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1013_ (.A1(_0340_),
    .A2(_0355_),
    .B(_0102_),
    .ZN(_0356_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1014_ (.A1(_0340_),
    .A2(_0355_),
    .B(_0356_),
    .ZN(_0357_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1015_ (.A1(_0329_),
    .A2(_0332_),
    .B(_0357_),
    .ZN(net41),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1016_ (.A1(_0106_),
    .A2(_0245_),
    .B(_0288_),
    .ZN(_0358_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1017_ (.A1(_0106_),
    .A2(_0247_),
    .B1(_0286_),
    .B2(_0093_),
    .C(_0358_),
    .ZN(_0359_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1018_ (.A1(_0189_),
    .A2(_0152_),
    .B(_0172_),
    .ZN(_0360_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1019_ (.A1(_0189_),
    .A2(_0156_),
    .B1(_0174_),
    .B2(_0169_),
    .C(_0360_),
    .ZN(_0361_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1020_ (.A1(\mprj.PS_R1_inst1.LUT_inst11.I1 ),
    .A2(_0119_),
    .B(_0130_),
    .ZN(_0362_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1021_ (.A1(_0239_),
    .A2(_0116_),
    .B1(_0132_),
    .B2(_0216_),
    .C(_0362_),
    .ZN(_0363_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1022_ (.A1(\mprj.PS_R1_inst1.LUT_inst13.I1 ),
    .A2(_0081_),
    .B(_0099_),
    .ZN(_0364_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1023_ (.A1(_0297_),
    .A2(_0076_),
    .B1(_0138_),
    .B2(\mprj.PS_R1_inst1.LUT_inst12.I1 ),
    .C(_0364_),
    .ZN(_0365_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1024_ (.A1(_0350_),
    .A2(_0363_),
    .A3(_0365_),
    .Z(_0366_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _1025_ (.A1(_0351_),
    .A2(_0361_),
    .A3(_0366_),
    .Z(_0367_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1026_ (.A1(_0146_),
    .A2(_0209_),
    .B(_0220_),
    .ZN(_0368_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1027_ (.A1(_0146_),
    .A2(_0205_),
    .B1(_0222_),
    .B2(_0126_),
    .C(_0368_),
    .ZN(_0369_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1028_ (.A1(_0352_),
    .A2(_0367_),
    .A3(_0369_),
    .Z(_0370_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1029_ (.A1(_0353_),
    .A2(_0359_),
    .A3(_0370_),
    .ZN(_0371_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1030_ (.A1(_0070_),
    .A2(_0319_),
    .ZN(_0372_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _1031_ (.I(\mprj.PS_Rx_inst7.LUT_inst1.i3 ),
    .ZN(_0373_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1032_ (.A1(_0373_),
    .A2(_0322_),
    .ZN(_0374_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1033_ (.A1(\mprj.PS_R1_inst1.LUT_inst2.I1 ),
    .A2(_0374_),
    .B(_0336_),
    .ZN(_0375_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1034_ (.A1(_0070_),
    .A2(_0334_),
    .B(_0372_),
    .C(_0375_),
    .ZN(_0376_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1035_ (.A1(_0354_),
    .A2(_0371_),
    .A3(_0376_),
    .Z(_0377_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1036_ (.A1(_0295_),
    .A2(\mprj.PS_Rx_inst8.LUT_inst1.i3 ),
    .ZN(_0378_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1037_ (.A1(_0295_),
    .A2(\mprj.PS_Rx_inst8.LUT_inst1.i3 ),
    .ZN(_0379_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1038_ (.A1(\mprj.PS_Rx_inst8.LUT_inst1.i4 ),
    .A2(_0379_),
    .ZN(_0380_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1039_ (.A1(_0378_),
    .A2(_0380_),
    .Z(_0381_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _1040_ (.I(_0381_),
    .Z(_0382_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1041_ (.A1(\mprj.PS_Rx_inst8.LUT_inst1.i3 ),
    .A2(\mprj.PS_Rx_inst8.LUT_inst1.i4 ),
    .Z(_0383_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1042_ (.A1(\mprj.PS_R1_inst1.LUT_inst1.i0 ),
    .A2(_0322_),
    .A3(_0383_),
    .Z(_0384_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _1043_ (.I(_0378_),
    .Z(_0385_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1044_ (.A1(_0078_),
    .A2(_0383_),
    .B(_0385_),
    .ZN(_0386_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1045_ (.A1(\mprj.PS_R1_inst1.LUT_inst1.i1 ),
    .A2(_0382_),
    .B1(_0384_),
    .B2(_0386_),
    .ZN(_0387_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1046_ (.A1(\mprj.PS_Rx_inst8.LUT_inst1.i4 ),
    .A2(_0377_),
    .A3(_0387_),
    .Z(_0388_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1047_ (.I(_0388_),
    .Z(\mprj.PS_Rx_inst8.carry_inst.O ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1048_ (.A1(_0103_),
    .A2(\mprj.PS_Rx_inst8.carry_inst.O ),
    .ZN(_0389_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _1049_ (.I(\mprj.PS_R1_inst1.LUT_inst15.I1 ),
    .ZN(_0390_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1050_ (.A1(net8),
    .A2(_0390_),
    .ZN(_0391_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _1051_ (.A1(\mprj.PS_Rx_inst8.LUT_inst1.i4 ),
    .A2(_0068_),
    .B1(_0391_),
    .B2(_0064_),
    .ZN(_0392_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1052_ (.A1(_0389_),
    .A2(_0392_),
    .ZN(net42),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1053_ (.A1(_0094_),
    .A2(_0316_),
    .B(_0333_),
    .ZN(_0393_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1054_ (.A1(_0094_),
    .A2(_0319_),
    .B1(_0336_),
    .B2(_0070_),
    .C(_0393_),
    .ZN(_0394_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1055_ (.A1(_0126_),
    .A2(_0249_),
    .B(_0289_),
    .ZN(_0395_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1056_ (.A1(_0127_),
    .A2(_0248_),
    .B1(_0287_),
    .B2(_0107_),
    .C(_0395_),
    .ZN(_0396_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1057_ (.A1(_0216_),
    .A2(_0152_),
    .B(_0173_),
    .ZN(_0397_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1058_ (.A1(_0216_),
    .A2(_0157_),
    .B1(_0175_),
    .B2(_0189_),
    .C(_0397_),
    .ZN(_0398_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1059_ (.A1(\mprj.PS_R1_inst1.LUT_inst12.I1 ),
    .A2(_0119_),
    .B(_0130_),
    .ZN(_0399_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1060_ (.A1(_0269_),
    .A2(_0116_),
    .B1(_0132_),
    .B2(\mprj.PS_R1_inst1.LUT_inst11.I1 ),
    .C(_0399_),
    .ZN(_0400_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1061_ (.A1(\mprj.PS_R1_inst1.LUT_inst14.I1 ),
    .A2(_0081_),
    .B(_0098_),
    .ZN(_0401_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1062_ (.A1(\mprj.PS_R1_inst1.LUT_inst14.I1 ),
    .A2(_0075_),
    .B1(_0138_),
    .B2(\mprj.PS_R1_inst1.LUT_inst13.I1 ),
    .C(_0401_),
    .ZN(_0402_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1063_ (.A1(_0365_),
    .A2(_0400_),
    .A3(_0402_),
    .ZN(_0403_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _1064_ (.A1(_0366_),
    .A2(_0398_),
    .A3(_0403_),
    .Z(_0404_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1065_ (.A1(_0169_),
    .A2(_0209_),
    .B(_0220_),
    .ZN(_0405_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1066_ (.A1(_0169_),
    .A2(_0205_),
    .B1(_0222_),
    .B2(_0146_),
    .C(_0405_),
    .ZN(_0406_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1067_ (.A1(_0367_),
    .A2(_0404_),
    .A3(_0406_),
    .Z(_0407_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1068_ (.A1(_0370_),
    .A2(_0396_),
    .A3(_0407_),
    .Z(_0408_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1069_ (.A1(_0371_),
    .A2(_0394_),
    .A3(_0408_),
    .Z(_0409_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1070_ (.A1(_0295_),
    .A2(\mprj.PS_Rx_inst8.LUT_inst1.i3 ),
    .B(\mprj.PS_Rx_inst8.LUT_inst1.i4 ),
    .ZN(_0410_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _1071_ (.I(_0410_),
    .Z(_0411_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1072_ (.A1(\mprj.PS_Rx_inst8.LUT_inst1.i4 ),
    .A2(_0379_),
    .ZN(_0412_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1073_ (.A1(_0378_),
    .A2(_0412_),
    .ZN(_0413_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1074_ (.A1(\mprj.PS_R1_inst1.LUT_inst1.i1 ),
    .A2(_0383_),
    .B(_0413_),
    .ZN(_0414_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1075_ (.A1(_0062_),
    .A2(_0381_),
    .ZN(_0415_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1076_ (.A1(_0062_),
    .A2(_0411_),
    .B(_0414_),
    .C(_0415_),
    .ZN(_0416_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _1077_ (.A1(_0409_),
    .A2(_0416_),
    .ZN(_0417_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1078_ (.A1(_0377_),
    .A2(_0417_),
    .Z(_0418_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1079_ (.A1(_0377_),
    .A2(_0417_),
    .B(_0103_),
    .ZN(_0419_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1080_ (.A1(_0060_),
    .A2(_0043_),
    .ZN(_0420_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _1081_ (.I(_0420_),
    .Z(_0421_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1082_ (.A1(_0418_),
    .A2(_0419_),
    .B(_0421_),
    .ZN(net43),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1083_ (.A1(_0107_),
    .A2(_0323_),
    .B(_0334_),
    .ZN(_0422_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1084_ (.A1(_0107_),
    .A2(_0320_),
    .B1(_0337_),
    .B2(_0094_),
    .C(_0422_),
    .ZN(_0423_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1085_ (.A1(\mprj.PS_R1_inst1.LUT_inst15.I1 ),
    .A2(_0080_),
    .B(_0098_),
    .ZN(_0424_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1086_ (.A1(\mprj.PS_R1_inst1.LUT_inst15.I1 ),
    .A2(_0075_),
    .B1(_0138_),
    .B2(\mprj.PS_R1_inst1.LUT_inst14.I1 ),
    .C(_0424_),
    .ZN(_0425_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1087_ (.A1(_0046_),
    .A2(_0425_),
    .Z(_0426_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1088_ (.A1(\mprj.PS_R1_inst1.LUT_inst13.I1 ),
    .A2(_0119_),
    .B(_0130_),
    .ZN(_0427_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1089_ (.A1(\mprj.PS_R1_inst1.LUT_inst13.I1 ),
    .A2(_0115_),
    .B1(_0132_),
    .B2(\mprj.PS_R1_inst1.LUT_inst12.I1 ),
    .C(_0427_),
    .ZN(_0428_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1090_ (.A1(_0402_),
    .A2(_0428_),
    .Z(_0429_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1091_ (.A1(_0426_),
    .A2(_0429_),
    .Z(_0430_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1092_ (.A1(_0239_),
    .A2(_0152_),
    .B(_0173_),
    .ZN(_0431_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1093_ (.A1(_0239_),
    .A2(_0157_),
    .B1(_0175_),
    .B2(_0216_),
    .C(_0431_),
    .ZN(_0432_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1094_ (.A1(_0403_),
    .A2(_0430_),
    .A3(_0432_),
    .ZN(_0433_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1095_ (.A1(_0189_),
    .A2(_0209_),
    .B(_0220_),
    .ZN(_0434_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1096_ (.A1(_0189_),
    .A2(_0205_),
    .B1(_0222_),
    .B2(_0169_),
    .C(_0434_),
    .ZN(_0435_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1097_ (.A1(_0433_),
    .A2(_0435_),
    .Z(_0436_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1098_ (.A1(_0147_),
    .A2(_0249_),
    .B(_0289_),
    .ZN(_0437_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1099_ (.A1(_0147_),
    .A2(_0248_),
    .B1(_0287_),
    .B2(_0127_),
    .C(_0437_),
    .ZN(_0438_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1100_ (.A1(_0367_),
    .A2(_0406_),
    .A3(_0438_),
    .ZN(_0439_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1101_ (.A1(_0436_),
    .A2(_0439_),
    .Z(_0440_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1102_ (.A1(_0408_),
    .A2(_0423_),
    .A3(_0440_),
    .Z(_0441_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1103_ (.A1(_0071_),
    .A2(_0382_),
    .ZN(_0442_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _1104_ (.I(_0413_),
    .Z(_0443_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1105_ (.A1(_0062_),
    .A2(_0383_),
    .B(_0443_),
    .ZN(_0444_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1106_ (.A1(_0071_),
    .A2(_0411_),
    .B(_0442_),
    .C(_0444_),
    .ZN(_0445_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1107_ (.A1(_0409_),
    .A2(_0441_),
    .A3(_0445_),
    .Z(_0446_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1108_ (.A1(_0051_),
    .A2(_0446_),
    .ZN(net44),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1109_ (.A1(_0127_),
    .A2(_0323_),
    .B(_0334_),
    .ZN(_0447_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1110_ (.A1(_0127_),
    .A2(_0320_),
    .B1(_0337_),
    .B2(_0107_),
    .C(_0447_),
    .ZN(_0448_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _1111_ (.I(\mprj.PS_R1_inst1.LUT_inst15.I1 ),
    .Z(_0449_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1112_ (.A1(_0136_),
    .A2(_0449_),
    .ZN(_0450_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _1113_ (.I(\mprj.PS_R1_inst1.LUT_inst14.I1 ),
    .ZN(_0451_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1114_ (.A1(_0052_),
    .A2(_0065_),
    .A3(_0451_),
    .ZN(_0452_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1115_ (.A1(_0046_),
    .A2(_0390_),
    .B(_0067_),
    .ZN(_0453_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1116_ (.A1(_0073_),
    .A2(_0450_),
    .B1(_0452_),
    .B2(_0453_),
    .ZN(_0454_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1117_ (.A1(\mprj.PS_R1_inst1.LUT_inst14.I1 ),
    .A2(_0119_),
    .B(_0130_),
    .ZN(_0455_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1118_ (.A1(\mprj.PS_R1_inst1.LUT_inst14.I1 ),
    .A2(_0116_),
    .B1(_0132_),
    .B2(_0297_),
    .C(_0455_),
    .ZN(_0456_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1119_ (.A1(_0454_),
    .A2(_0456_),
    .Z(_0457_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1120_ (.A1(_0269_),
    .A2(_0152_),
    .B(_0173_),
    .ZN(_0458_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1121_ (.A1(_0269_),
    .A2(_0157_),
    .B1(_0175_),
    .B2(_0239_),
    .C(_0458_),
    .ZN(_0459_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1122_ (.A1(_0429_),
    .A2(_0457_),
    .A3(_0459_),
    .Z(_0460_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1123_ (.A1(_0216_),
    .A2(_0209_),
    .B(_0220_),
    .ZN(_0461_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1124_ (.A1(_0216_),
    .A2(_0205_),
    .B1(_0222_),
    .B2(_0189_),
    .C(_0461_),
    .ZN(_0462_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1125_ (.A1(_0433_),
    .A2(_0460_),
    .A3(_0462_),
    .Z(_0463_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1126_ (.A1(_0169_),
    .A2(_0245_),
    .B(_0288_),
    .ZN(_0464_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1127_ (.A1(_0170_),
    .A2(_0247_),
    .B1(_0286_),
    .B2(_0146_),
    .C(_0464_),
    .ZN(_0465_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1128_ (.A1(_0404_),
    .A2(_0465_),
    .Z(_0466_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1129_ (.A1(_0436_),
    .A2(_0463_),
    .A3(_0466_),
    .Z(_0467_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _1130_ (.A1(_0440_),
    .A2(_0448_),
    .A3(_0467_),
    .Z(_0468_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1131_ (.A1(_0094_),
    .A2(_0385_),
    .B(_0411_),
    .ZN(_0469_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1132_ (.A1(_0094_),
    .A2(_0382_),
    .B1(_0443_),
    .B2(_0071_),
    .C(_0469_),
    .ZN(_0470_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1133_ (.A1(_0441_),
    .A2(_0470_),
    .Z(_0471_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1134_ (.A1(_0468_),
    .A2(_0471_),
    .Z(_0472_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1135_ (.A1(_0468_),
    .A2(_0471_),
    .B(_0103_),
    .ZN(_0473_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1136_ (.A1(_0472_),
    .A2(_0473_),
    .B(_0421_),
    .ZN(net45),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1137_ (.A1(_0107_),
    .A2(_0385_),
    .B(_0411_),
    .ZN(_0474_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1138_ (.A1(_0107_),
    .A2(_0382_),
    .B1(_0443_),
    .B2(_0094_),
    .C(_0474_),
    .ZN(_0475_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1139_ (.A1(_0147_),
    .A2(_0323_),
    .B(_0334_),
    .ZN(_0476_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1140_ (.A1(_0147_),
    .A2(_0320_),
    .B1(_0337_),
    .B2(_0127_),
    .C(_0476_),
    .ZN(_0477_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1141_ (.A1(_0189_),
    .A2(_0249_),
    .B(_0289_),
    .ZN(_0478_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1142_ (.A1(_0190_),
    .A2(_0248_),
    .B1(_0287_),
    .B2(_0170_),
    .C(_0478_),
    .ZN(_0479_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1143_ (.A1(_0297_),
    .A2(_0151_),
    .B(_0172_),
    .ZN(_0480_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1144_ (.A1(_0297_),
    .A2(_0156_),
    .B1(_0174_),
    .B2(_0269_),
    .C(_0480_),
    .ZN(_0481_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1145_ (.A1(_0426_),
    .A2(_0481_),
    .Z(_0482_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1146_ (.A1(\mprj.PS_R1_inst1.LUT_inst14.I1 ),
    .A2(_0117_),
    .Z(_0483_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1147_ (.A1(_0449_),
    .A2(_0130_),
    .ZN(_0484_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1148_ (.A1(_0449_),
    .A2(_0116_),
    .B1(_0132_),
    .B2(_0483_),
    .C(_0484_),
    .ZN(_0485_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1149_ (.A1(_0086_),
    .A2(_0454_),
    .A3(_0485_),
    .Z(_0486_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1150_ (.A1(_0457_),
    .A2(_0482_),
    .A3(_0486_),
    .Z(_0487_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1151_ (.A1(_0239_),
    .A2(_0209_),
    .B(_0220_),
    .ZN(_0488_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1152_ (.A1(_0239_),
    .A2(_0205_),
    .B1(_0222_),
    .B2(_0216_),
    .C(_0488_),
    .ZN(_0489_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1153_ (.A1(_0460_),
    .A2(_0487_),
    .A3(_0489_),
    .ZN(_0490_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1154_ (.A1(_0463_),
    .A2(_0479_),
    .A3(_0490_),
    .ZN(_0491_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1155_ (.A1(_0467_),
    .A2(_0477_),
    .A3(_0491_),
    .Z(_0492_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1156_ (.A1(_0475_),
    .A2(_0492_),
    .Z(_0493_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1157_ (.A1(_0468_),
    .A2(_0493_),
    .Z(_0494_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1158_ (.A1(_0468_),
    .A2(_0493_),
    .B(_0103_),
    .ZN(_0495_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1159_ (.A1(_0494_),
    .A2(_0495_),
    .B(_0421_),
    .ZN(net46),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1160_ (.A1(_0170_),
    .A2(_0323_),
    .B(_0333_),
    .ZN(_0496_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1161_ (.A1(_0170_),
    .A2(_0319_),
    .B1(_0337_),
    .B2(_0147_),
    .C(_0496_),
    .ZN(_0497_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1162_ (.A1(_0216_),
    .A2(_0249_),
    .B(_0288_),
    .ZN(_0498_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1163_ (.A1(_0217_),
    .A2(_0247_),
    .B1(_0286_),
    .B2(_0190_),
    .C(_0498_),
    .ZN(_0499_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1164_ (.A1(_0330_),
    .A2(_0152_),
    .B(_0173_),
    .ZN(_0500_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1165_ (.A1(_0330_),
    .A2(_0157_),
    .B1(_0175_),
    .B2(_0297_),
    .C(_0500_),
    .ZN(_0501_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1166_ (.A1(_0486_),
    .A2(_0501_),
    .Z(_0502_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1167_ (.A1(_0136_),
    .A2(\mprj.PS_Rx_inst3.LUT_inst1.i3 ),
    .A3(_0451_),
    .ZN(_0503_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1168_ (.A1(_0104_),
    .A2(_0450_),
    .ZN(_0504_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1169_ (.A1(_0112_),
    .A2(_0449_),
    .A3(_0114_),
    .ZN(_0505_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1170_ (.A1(_0503_),
    .A2(_0504_),
    .B(_0505_),
    .ZN(_0506_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1171_ (.A1(_0269_),
    .A2(_0209_),
    .B(_0219_),
    .ZN(_0507_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1172_ (.A1(_0269_),
    .A2(_0204_),
    .B1(_0221_),
    .B2(_0239_),
    .C(_0507_),
    .ZN(_0508_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1173_ (.A1(_0506_),
    .A2(_0508_),
    .Z(_0509_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1174_ (.A1(_0487_),
    .A2(_0502_),
    .A3(_0509_),
    .Z(_0510_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1175_ (.A1(_0490_),
    .A2(_0499_),
    .A3(_0510_),
    .ZN(_0511_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _1176_ (.A1(_0491_),
    .A2(_0497_),
    .A3(_0511_),
    .Z(_0512_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1177_ (.A1(_0127_),
    .A2(_0385_),
    .B(_0411_),
    .ZN(_0513_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1178_ (.A1(_0127_),
    .A2(_0382_),
    .B1(_0443_),
    .B2(_0107_),
    .C(_0513_),
    .ZN(_0514_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1179_ (.A1(_0492_),
    .A2(_0512_),
    .A3(_0514_),
    .Z(_0515_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1180_ (.A1(_0051_),
    .A2(_0515_),
    .ZN(net48),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1181_ (.A1(_0147_),
    .A2(_0385_),
    .B(_0411_),
    .ZN(_0516_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1182_ (.A1(_0147_),
    .A2(_0382_),
    .B1(_0443_),
    .B2(_0127_),
    .C(_0516_),
    .ZN(_0517_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1183_ (.A1(_0297_),
    .A2(_0209_),
    .B(_0220_),
    .ZN(_0518_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1184_ (.A1(_0297_),
    .A2(_0204_),
    .B1(_0222_),
    .B2(_0269_),
    .C(_0518_),
    .ZN(_0519_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1185_ (.A1(_0330_),
    .A2(_0149_),
    .B(_0175_),
    .ZN(_0520_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1186_ (.A1(_0449_),
    .A2(_0157_),
    .ZN(_0521_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1187_ (.A1(_0449_),
    .A2(_0173_),
    .B(_0520_),
    .C(_0521_),
    .ZN(_0522_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1188_ (.A1(_0055_),
    .A2(_0522_),
    .Z(_0523_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1189_ (.A1(_0502_),
    .A2(_0519_),
    .A3(_0523_),
    .Z(_0524_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1190_ (.A1(_0239_),
    .A2(_0249_),
    .B(_0289_),
    .ZN(_0525_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1191_ (.A1(_0240_),
    .A2(_0248_),
    .B1(_0287_),
    .B2(_0217_),
    .C(_0525_),
    .ZN(_0526_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1192_ (.A1(_0510_),
    .A2(_0524_),
    .A3(_0526_),
    .Z(_0527_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1193_ (.A1(_0190_),
    .A2(_0323_),
    .B(_0334_),
    .ZN(_0528_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1194_ (.A1(_0190_),
    .A2(_0320_),
    .B1(_0337_),
    .B2(_0170_),
    .C(_0528_),
    .ZN(_0529_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1195_ (.A1(_0511_),
    .A2(_0527_),
    .A3(_0529_),
    .Z(_0530_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _1196_ (.A1(_0517_),
    .A2(_0530_),
    .ZN(_0531_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1197_ (.A1(_0512_),
    .A2(_0531_),
    .ZN(_0532_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1198_ (.A1(_0512_),
    .A2(_0531_),
    .Z(_0533_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _1199_ (.A1(_0051_),
    .A2(_0532_),
    .A3(_0533_),
    .B(_0420_),
    .ZN(net49),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1200_ (.A1(_0217_),
    .A2(_0316_),
    .B(_0333_),
    .ZN(_0534_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1201_ (.A1(_0217_),
    .A2(_0319_),
    .B1(_0336_),
    .B2(_0190_),
    .C(_0534_),
    .ZN(_0535_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1202_ (.A1(_0269_),
    .A2(_0249_),
    .B(_0289_),
    .ZN(_0536_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1203_ (.A1(_0270_),
    .A2(_0248_),
    .B1(_0287_),
    .B2(_0240_),
    .C(_0536_),
    .ZN(_0537_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1204_ (.A1(_0330_),
    .A2(_0208_),
    .B(_0219_),
    .ZN(_0538_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1205_ (.A1(_0330_),
    .A2(_0204_),
    .B1(_0221_),
    .B2(_0297_),
    .C(_0538_),
    .ZN(_0539_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1206_ (.A1(_0144_),
    .A2(_0390_),
    .ZN(_0540_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1207_ (.A1(_0112_),
    .A2(\mprj.PS_Rx_inst4.LUT_inst1.i3 ),
    .ZN(_0541_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1208_ (.A1(_0112_),
    .A2(_0449_),
    .B1(_0541_),
    .B2(_0330_),
    .C(_0154_),
    .ZN(_0542_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1209_ (.A1(_0155_),
    .A2(_0540_),
    .B(_0542_),
    .ZN(_0543_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1210_ (.A1(_0506_),
    .A2(_0539_),
    .A3(_0543_),
    .Z(_0544_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1211_ (.A1(_0523_),
    .A2(_0544_),
    .Z(_0545_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1212_ (.A1(_0524_),
    .A2(_0537_),
    .A3(_0545_),
    .Z(_0546_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_4 _1213_ (.A1(_0527_),
    .A2(_0535_),
    .A3(_0546_),
    .ZN(_0547_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1214_ (.A1(_0170_),
    .A2(_0385_),
    .B(_0411_),
    .ZN(_0548_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1215_ (.A1(_0170_),
    .A2(_0382_),
    .B1(_0443_),
    .B2(_0147_),
    .C(_0548_),
    .ZN(_0549_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1216_ (.A1(_0530_),
    .A2(_0547_),
    .A3(_0549_),
    .Z(_0550_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1217_ (.A1(_0051_),
    .A2(_0550_),
    .ZN(net50),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1218_ (.A1(_0190_),
    .A2(_0385_),
    .B(_0411_),
    .ZN(_0551_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1219_ (.A1(_0190_),
    .A2(_0382_),
    .B1(_0443_),
    .B2(_0170_),
    .C(_0551_),
    .ZN(_0552_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1220_ (.A1(_0240_),
    .A2(_0323_),
    .B(_0333_),
    .ZN(_0553_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1221_ (.A1(_0240_),
    .A2(_0319_),
    .B1(_0336_),
    .B2(_0217_),
    .C(_0553_),
    .ZN(_0554_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1222_ (.A1(_0297_),
    .A2(_0249_),
    .B(_0289_),
    .ZN(_0555_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1223_ (.A1(_0298_),
    .A2(_0248_),
    .B1(_0287_),
    .B2(_0270_),
    .C(_0555_),
    .ZN(_0556_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1224_ (.A1(_0449_),
    .A2(_0205_),
    .ZN(_0557_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1225_ (.A1(_0330_),
    .A2(_0206_),
    .B(_0222_),
    .ZN(_0558_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1226_ (.A1(_0449_),
    .A2(_0220_),
    .B(_0557_),
    .C(_0558_),
    .ZN(_0559_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1227_ (.A1(_0055_),
    .A2(_0543_),
    .A3(_0559_),
    .Z(_0560_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1228_ (.A1(_0545_),
    .A2(_0556_),
    .A3(_0560_),
    .ZN(_0561_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _1229_ (.A1(_0546_),
    .A2(_0554_),
    .A3(_0561_),
    .Z(_0562_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1230_ (.A1(_0552_),
    .A2(_0562_),
    .Z(_0563_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1231_ (.A1(_0547_),
    .A2(_0563_),
    .B(_0051_),
    .ZN(_0564_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1232_ (.A1(_0547_),
    .A2(_0563_),
    .B(_0564_),
    .ZN(_0565_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1233_ (.A1(_0421_),
    .A2(_0565_),
    .ZN(net51),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1234_ (.A1(_0217_),
    .A2(_0385_),
    .B(_0411_),
    .ZN(_0566_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1235_ (.A1(_0217_),
    .A2(_0382_),
    .B1(_0443_),
    .B2(_0190_),
    .C(_0566_),
    .ZN(_0567_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1236_ (.A1(_0270_),
    .A2(_0323_),
    .B(_0334_),
    .ZN(_0568_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1237_ (.A1(_0270_),
    .A2(_0320_),
    .B1(_0337_),
    .B2(_0240_),
    .C(_0568_),
    .ZN(_0569_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1238_ (.A1(_0154_),
    .A2(\mprj.PS_Rx_inst5.LUT_inst1.i3 ),
    .A3(_0451_),
    .ZN(_0570_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1239_ (.A1(_0144_),
    .A2(_0390_),
    .B(_0187_),
    .ZN(_0571_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1240_ (.A1(_0390_),
    .A2(_0203_),
    .B1(_0570_),
    .B2(_0571_),
    .ZN(_0572_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1241_ (.A1(_0330_),
    .A2(_0249_),
    .B(_0289_),
    .ZN(_0573_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1242_ (.A1(_0330_),
    .A2(_0248_),
    .B1(_0287_),
    .B2(_0298_),
    .C(_0573_),
    .ZN(_0574_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1243_ (.A1(_0560_),
    .A2(_0572_),
    .A3(_0574_),
    .Z(_0575_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _1244_ (.A1(_0561_),
    .A2(_0569_),
    .A3(_0575_),
    .Z(_0576_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_4 _1245_ (.A1(_0567_),
    .A2(_0576_),
    .ZN(_0577_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1246_ (.A1(_0562_),
    .A2(_0577_),
    .B(_0103_),
    .ZN(_0578_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1247_ (.A1(_0562_),
    .A2(_0577_),
    .B(_0578_),
    .ZN(net52),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1248_ (.A1(_0240_),
    .A2(_0385_),
    .B(_0410_),
    .ZN(_0579_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1249_ (.A1(_0240_),
    .A2(_0381_),
    .B1(_0443_),
    .B2(_0217_),
    .C(_0579_),
    .ZN(_0580_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1250_ (.A1(_0298_),
    .A2(_0323_),
    .B(_0334_),
    .ZN(_0581_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1251_ (.A1(_0298_),
    .A2(_0320_),
    .B1(_0337_),
    .B2(_0270_),
    .C(_0581_),
    .ZN(_0582_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1252_ (.A1(_0237_),
    .A2(_0390_),
    .A3(_0244_),
    .ZN(_0583_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1253_ (.A1(_0249_),
    .A2(_0583_),
    .ZN(_0584_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1254_ (.A1(_0451_),
    .A2(_0243_),
    .ZN(_0585_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _1255_ (.I(_0449_),
    .Z(_0586_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1256_ (.A1(_0586_),
    .A2(_0289_),
    .ZN(_0587_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1257_ (.A1(_0287_),
    .A2(_0585_),
    .B(_0587_),
    .ZN(_0588_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1258_ (.A1(_0584_),
    .A2(_0588_),
    .ZN(_0589_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1259_ (.A1(_0086_),
    .A2(_0572_),
    .A3(_0589_),
    .Z(_0590_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _1260_ (.A1(_0575_),
    .A2(_0582_),
    .A3(_0590_),
    .Z(_0591_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1261_ (.A1(_0580_),
    .A2(_0591_),
    .Z(_0592_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1262_ (.A1(_0576_),
    .A2(_0592_),
    .B(_0050_),
    .ZN(_0593_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1263_ (.A1(_0576_),
    .A2(_0592_),
    .B(_0593_),
    .ZN(_0594_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1264_ (.A1(_0421_),
    .A2(_0594_),
    .ZN(net53),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1265_ (.A1(_0331_),
    .A2(_0323_),
    .B(_0334_),
    .ZN(_0595_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1266_ (.A1(_0331_),
    .A2(_0320_),
    .B1(_0337_),
    .B2(_0298_),
    .C(_0595_),
    .ZN(_0596_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1267_ (.A1(_0590_),
    .A2(_0596_),
    .Z(_0597_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1268_ (.A1(_0270_),
    .A2(_0378_),
    .B(_0410_),
    .ZN(_0598_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1269_ (.A1(_0270_),
    .A2(_0381_),
    .B1(_0413_),
    .B2(_0240_),
    .C(_0598_),
    .ZN(_0599_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _1270_ (.I(\mprj.PS_Rx_inst6.LUT_inst1.i3 ),
    .ZN(_0600_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1271_ (.A1(_0187_),
    .A2(_0600_),
    .A3(_0331_),
    .ZN(_0601_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1272_ (.A1(_0201_),
    .A2(_0586_),
    .B(_0242_),
    .ZN(_0602_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1273_ (.A1(_0601_),
    .A2(_0602_),
    .B(_0583_),
    .ZN(_0603_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_4 _1274_ (.A1(_0597_),
    .A2(_0599_),
    .A3(_0603_),
    .Z(_0604_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1275_ (.A1(_0591_),
    .A2(_0604_),
    .Z(_0605_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1276_ (.A1(_0591_),
    .A2(_0604_),
    .B(_0103_),
    .ZN(_0606_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1277_ (.A1(_0605_),
    .A2(_0606_),
    .B(_0421_),
    .ZN(net54),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1278_ (.A1(_0298_),
    .A2(_0385_),
    .B(_0410_),
    .ZN(_0607_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1279_ (.A1(_0298_),
    .A2(_0381_),
    .B1(_0413_),
    .B2(_0270_),
    .C(_0607_),
    .ZN(_0608_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1280_ (.A1(_0586_),
    .A2(_0320_),
    .ZN(_0609_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1281_ (.A1(_0331_),
    .A2(_0374_),
    .B(_0337_),
    .ZN(_0610_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1282_ (.A1(_0586_),
    .A2(_0334_),
    .B(_0609_),
    .C(_0610_),
    .ZN(_0611_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1283_ (.A1(_0055_),
    .A2(_0611_),
    .Z(_0612_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1284_ (.A1(_0608_),
    .A2(_0612_),
    .Z(_0613_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1285_ (.A1(_0597_),
    .A2(_0613_),
    .B(_0050_),
    .ZN(_0614_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1286_ (.A1(_0597_),
    .A2(_0613_),
    .B(_0614_),
    .ZN(_0615_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1287_ (.A1(_0421_),
    .A2(_0615_),
    .ZN(net55),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1288_ (.A1(_0331_),
    .A2(_0378_),
    .B(_0410_),
    .ZN(_0616_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1289_ (.A1(_0331_),
    .A2(_0381_),
    .B1(_0413_),
    .B2(_0298_),
    .C(_0616_),
    .ZN(_0617_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1290_ (.A1(_0237_),
    .A2(_0373_),
    .A3(_0331_),
    .ZN(_0618_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1291_ (.A1(_0242_),
    .A2(_0586_),
    .B(_0322_),
    .ZN(_0619_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1292_ (.A1(_0586_),
    .A2(_0318_),
    .B1(_0618_),
    .B2(_0619_),
    .ZN(_0620_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1293_ (.A1(_0603_),
    .A2(_0620_),
    .Z(_0621_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1294_ (.A1(_0617_),
    .A2(_0621_),
    .Z(_0622_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1295_ (.A1(_0612_),
    .A2(_0622_),
    .B(_0050_),
    .ZN(_0623_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1296_ (.A1(_0612_),
    .A2(_0622_),
    .B(_0623_),
    .ZN(_0624_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1297_ (.A1(_0421_),
    .A2(_0624_),
    .ZN(net56),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1298_ (.A1(_0331_),
    .A2(_0383_),
    .B(_0443_),
    .ZN(_0625_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1299_ (.A1(_0586_),
    .A2(_0382_),
    .ZN(_0626_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1300_ (.A1(_0586_),
    .A2(_0411_),
    .B(_0625_),
    .C(_0626_),
    .ZN(_0627_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1301_ (.A1(_0086_),
    .A2(_0620_),
    .Z(_0628_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1302_ (.A1(_0627_),
    .A2(_0628_),
    .B(_0051_),
    .ZN(_0629_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1303_ (.A1(_0627_),
    .A2(_0628_),
    .B(_0629_),
    .ZN(_0630_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1304_ (.I(_0630_),
    .ZN(net57),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1305_ (.A1(_0322_),
    .A2(\mprj.PS_Rx_inst8.LUT_inst1.i3 ),
    .ZN(_0631_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1306_ (.A1(_0322_),
    .A2(_0586_),
    .B1(_0631_),
    .B2(_0331_),
    .ZN(_0632_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1307_ (.A1(_0586_),
    .A2(_0380_),
    .B1(_0632_),
    .B2(\mprj.PS_Rx_inst8.LUT_inst1.i4 ),
    .C(_0050_),
    .ZN(_0633_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1308_ (.I(_0633_),
    .ZN(_0634_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1309_ (.A1(_0421_),
    .A2(_0634_),
    .ZN(net59),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1310_ (.A1(_0051_),
    .A2(_0055_),
    .B(_0421_),
    .ZN(net60),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1311_ (.I(net1),
    .ZN(net34),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1312_ (.A1(net4),
    .A2(net2),
    .A3(_0034_),
    .ZN(_0635_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1313_ (.A1(_0039_),
    .A2(_0635_),
    .ZN(_0636_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 _1314_ (.I(_0636_),
    .Z(_0637_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1315_ (.A1(net14),
    .A2(_0637_),
    .ZN(_0638_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1316_ (.A1(_0035_),
    .A2(_0637_),
    .B(_0638_),
    .ZN(_0000_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1317_ (.A1(net21),
    .A2(_0637_),
    .ZN(_0639_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1318_ (.A1(_0053_),
    .A2(_0637_),
    .B(_0639_),
    .ZN(_0001_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1319_ (.I0(net22),
    .I1(_0063_),
    .S(_0637_),
    .Z(_0640_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1320_ (.I(_0640_),
    .Z(_0002_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1321_ (.I0(net23),
    .I1(_0071_),
    .S(_0637_),
    .Z(_0641_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1322_ (.I(_0641_),
    .Z(_0003_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _1323_ (.I(_0636_),
    .Z(_0642_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1324_ (.I0(net24),
    .I1(_0094_),
    .S(_0642_),
    .Z(_0643_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1325_ (.I(_0643_),
    .Z(_0004_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1326_ (.I0(net25),
    .I1(_0107_),
    .S(_0642_),
    .Z(_0644_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1327_ (.I(_0644_),
    .Z(_0005_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1328_ (.I0(net26),
    .I1(_0127_),
    .S(_0642_),
    .Z(_0645_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1329_ (.I(_0645_),
    .Z(_0006_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1330_ (.I0(net27),
    .I1(_0147_),
    .S(_0642_),
    .Z(_0646_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1331_ (.I(_0646_),
    .Z(_0007_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1332_ (.I0(net28),
    .I1(_0170_),
    .S(_0642_),
    .Z(_0647_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1333_ (.I(_0647_),
    .Z(_0008_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1334_ (.I0(net29),
    .I1(_0190_),
    .S(_0642_),
    .Z(_0648_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1335_ (.I(_0648_),
    .Z(_0009_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1336_ (.I0(net15),
    .I1(_0217_),
    .S(_0642_),
    .Z(_0649_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1337_ (.I(_0649_),
    .Z(_0010_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1338_ (.I0(net16),
    .I1(_0240_),
    .S(_0642_),
    .Z(_0650_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1339_ (.I(_0650_),
    .Z(_0011_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1340_ (.I0(net17),
    .I1(_0270_),
    .S(_0642_),
    .Z(_0651_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1341_ (.I(_0651_),
    .Z(_0012_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1342_ (.I0(net18),
    .I1(_0298_),
    .S(_0642_),
    .Z(_0652_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1343_ (.I(_0652_),
    .Z(_0013_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1344_ (.A1(net19),
    .A2(_0637_),
    .ZN(_0653_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1345_ (.A1(_0451_),
    .A2(_0637_),
    .B(_0653_),
    .ZN(_0014_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1346_ (.A1(net20),
    .A2(_0637_),
    .ZN(_0654_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1347_ (.A1(_0390_),
    .A2(_0637_),
    .B(_0654_),
    .ZN(_0015_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1348_ (.A1(_0042_),
    .A2(_0635_),
    .ZN(_0655_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _1349_ (.I(_0655_),
    .Z(_0656_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _1350_ (.I(_0655_),
    .Z(_0657_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1351_ (.A1(net14),
    .A2(_0657_),
    .ZN(_0658_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1352_ (.A1(_0047_),
    .A2(_0656_),
    .B(_0658_),
    .ZN(_0016_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1353_ (.A1(net21),
    .A2(_0657_),
    .ZN(_0659_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1354_ (.A1(_0052_),
    .A2(_0656_),
    .B(_0659_),
    .ZN(_0017_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1355_ (.I0(net22),
    .I1(_0065_),
    .S(_0655_),
    .Z(_0660_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1356_ (.I(_0660_),
    .Z(_0018_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1357_ (.A1(net23),
    .A2(_0657_),
    .ZN(_0661_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1358_ (.A1(_0136_),
    .A2(_0656_),
    .B(_0661_),
    .ZN(_0019_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1359_ (.I0(net24),
    .I1(\mprj.PS_Rx_inst3.LUT_inst1.i3 ),
    .S(_0655_),
    .Z(_0662_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1360_ (.I(_0662_),
    .Z(_0020_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1361_ (.A1(net25),
    .A2(_0657_),
    .ZN(_0663_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1362_ (.A1(_0112_),
    .A2(_0656_),
    .B(_0663_),
    .ZN(_0021_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1363_ (.I0(net26),
    .I1(\mprj.PS_Rx_inst4.LUT_inst1.i3 ),
    .S(_0655_),
    .Z(_0664_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1364_ (.I(_0664_),
    .Z(_0022_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1365_ (.A1(net27),
    .A2(_0657_),
    .ZN(_0665_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1366_ (.A1(_0154_),
    .A2(_0656_),
    .B(_0665_),
    .ZN(_0023_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1367_ (.I0(net28),
    .I1(\mprj.PS_Rx_inst5.LUT_inst1.i3 ),
    .S(_0655_),
    .Z(_0666_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1368_ (.I(_0666_),
    .Z(_0024_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1369_ (.A1(net29),
    .A2(_0657_),
    .ZN(_0667_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1370_ (.A1(_0201_),
    .A2(_0656_),
    .B(_0667_),
    .ZN(_0025_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1371_ (.A1(net15),
    .A2(_0657_),
    .ZN(_0668_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1372_ (.A1(_0600_),
    .A2(_0656_),
    .B(_0668_),
    .ZN(_0026_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1373_ (.A1(net16),
    .A2(_0657_),
    .ZN(_0669_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1374_ (.A1(_0242_),
    .A2(_0656_),
    .B(_0669_),
    .ZN(_0027_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1375_ (.A1(net17),
    .A2(_0657_),
    .ZN(_0670_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1376_ (.A1(_0373_),
    .A2(_0656_),
    .B(_0670_),
    .ZN(_0028_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1377_ (.A1(net18),
    .A2(_0657_),
    .ZN(_0671_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1378_ (.A1(_0322_),
    .A2(_0656_),
    .B(_0671_),
    .ZN(_0029_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1379_ (.I0(net19),
    .I1(\mprj.PS_Rx_inst8.LUT_inst1.i3 ),
    .S(_0655_),
    .Z(_0672_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1380_ (.I(_0672_),
    .Z(_0030_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1381_ (.I0(net20),
    .I1(\mprj.PS_Rx_inst8.LUT_inst1.i4 ),
    .S(_0655_),
    .Z(_0673_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1382_ (.I(_0673_),
    .Z(_0031_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1383_ (.D(\mprj.PS_R1_inst1.LUT_inst1.i0 ),
    .CLK(net71),
    .Q(net32),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1384_ (.D(\mprj.PS_Rx_inst8.carry_inst.O ),
    .CLK(net68),
    .Q(net33),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1385_ (.D(_0000_),
    .CLK(net71),
    .Q(\mprj.PS_R1_inst1.LUT_inst1.i0 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1386_ (.D(_0001_),
    .CLK(net70),
    .Q(\mprj.PS_R1_inst1.LUT_inst1.i1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1387_ (.D(_0002_),
    .CLK(net70),
    .Q(\mprj.PS_R1_inst1.LUT_inst2.I1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1388_ (.D(_0003_),
    .CLK(net68),
    .Q(\mprj.PS_R1_inst1.LUT_inst3.I1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1389_ (.D(_0004_),
    .CLK(net70),
    .Q(\mprj.PS_R1_inst1.LUT_inst4.I1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1390_ (.D(_0005_),
    .CLK(net70),
    .Q(\mprj.PS_R1_inst1.LUT_inst5.I1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1391_ (.D(_0006_),
    .CLK(net68),
    .Q(\mprj.PS_R1_inst1.LUT_inst6.I1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1392_ (.D(_0007_),
    .CLK(net68),
    .Q(\mprj.PS_R1_inst1.LUT_inst7.I1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1393_ (.D(_0008_),
    .CLK(net69),
    .Q(\mprj.PS_R1_inst1.LUT_inst8.I1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1394_ (.D(_0009_),
    .CLK(net69),
    .Q(\mprj.PS_R1_inst1.LUT_inst10.I0 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1395_ (.D(_0010_),
    .CLK(net69),
    .Q(\mprj.PS_R1_inst1.LUT_inst10.I1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1396_ (.D(_0011_),
    .CLK(net71),
    .Q(\mprj.PS_R1_inst1.LUT_inst11.I1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1397_ (.D(_0012_),
    .CLK(net71),
    .Q(\mprj.PS_R1_inst1.LUT_inst12.I1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1398_ (.D(_0013_),
    .CLK(net68),
    .Q(\mprj.PS_R1_inst1.LUT_inst13.I1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1399_ (.D(_0014_),
    .CLK(net71),
    .Q(\mprj.PS_R1_inst1.LUT_inst14.I1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1400_ (.D(_0015_),
    .CLK(net69),
    .Q(\mprj.PS_R1_inst1.LUT_inst15.I1 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1401_ (.D(_0016_),
    .CLK(net68),
    .Q(\mprj.PS_R1_inst1.LUT_inst1.i3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1402_ (.D(_0017_),
    .CLK(net70),
    .Q(\mprj.PS_R1_inst1.LUT_inst1.i4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1403_ (.D(_0018_),
    .CLK(net69),
    .Q(\mprj.PS_Rx_inst2.LUT_inst1.i3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1404_ (.D(_0019_),
    .CLK(net69),
    .Q(\mprj.PS_Rx_inst2.LUT_inst1.i4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1405_ (.D(_0020_),
    .CLK(net68),
    .Q(\mprj.PS_Rx_inst3.LUT_inst1.i3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1406_ (.D(_0021_),
    .CLK(net70),
    .Q(\mprj.PS_Rx_inst3.LUT_inst1.i4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1407_ (.D(_0022_),
    .CLK(net70),
    .Q(\mprj.PS_Rx_inst4.LUT_inst1.i3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1408_ (.D(_0023_),
    .CLK(net70),
    .Q(\mprj.PS_Rx_inst4.LUT_inst1.i4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1409_ (.D(_0024_),
    .CLK(net70),
    .Q(\mprj.PS_Rx_inst5.LUT_inst1.i3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1410_ (.D(_0025_),
    .CLK(net68),
    .Q(\mprj.PS_Rx_inst5.LUT_inst1.i4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1411_ (.D(_0026_),
    .CLK(net70),
    .Q(\mprj.PS_Rx_inst6.LUT_inst1.i3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1412_ (.D(_0027_),
    .CLK(net71),
    .Q(\mprj.PS_Rx_inst6.LUT_inst1.i4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1413_ (.D(_0028_),
    .CLK(net69),
    .Q(\mprj.PS_Rx_inst7.LUT_inst1.i3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1414_ (.D(_0029_),
    .CLK(net68),
    .Q(\mprj.PS_Rx_inst7.LUT_inst1.i4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1415_ (.D(_0030_),
    .CLK(net68),
    .Q(\mprj.PS_Rx_inst8.LUT_inst1.i3 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _1416_ (.D(_0031_),
    .CLK(net71),
    .Q(\mprj.PS_Rx_inst8.LUT_inst1.i4 ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_73 (.ZN(net73),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_74 (.ZN(net74),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_75 (.ZN(net75),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_76 (.ZN(net76),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_77 (.ZN(net77),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_78 (.ZN(net78),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_79 (.ZN(net79),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_80 (.ZN(net80),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_81 (.ZN(net81),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_82 (.ZN(net82),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_83 (.ZN(net83),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_84 (.ZN(net84),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_85 (.ZN(net85),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_86 (.ZN(net86),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_87 (.ZN(net87),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_88 (.ZN(net88),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_89 (.ZN(net89),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_90 (.ZN(net90),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_91 (.ZN(net91),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_92 (.ZN(net92),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_93 (.ZN(net93),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_94 (.ZN(net94),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_95 (.ZN(net95),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_96 (.ZN(net96),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_97 (.ZN(net97),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_98 (.ZN(net98),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_99 (.ZN(net99),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_100 (.ZN(net100),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_101 (.ZN(net101),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_102 (.ZN(net102),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_103 (.ZN(net103),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_104 (.ZN(net104),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_105 (.ZN(net105),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_106 (.ZN(net106),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_107 (.ZN(net107),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_108 (.ZN(net108),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_109 (.ZN(net109),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_110 (.ZN(net110),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_111 (.ZN(net111),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_112 (.ZN(net112),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_113 (.ZN(net113),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_114 (.ZN(net114),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_115 (.ZN(net115),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_116 (.ZN(net116),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_117 (.ZN(net117),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_118 (.ZN(net118),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_119 (.ZN(net119),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_120 (.ZN(net120),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_121 (.ZN(net121),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_122 (.ZN(net122),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_123 (.ZN(net123),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_124 (.ZN(net124),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_125 (.ZN(net125),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_126 (.ZN(net126),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_127 (.ZN(net127),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_128 (.ZN(net128),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_129 (.ZN(net129),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_130 (.ZN(net130),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_131 (.ZN(net131),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_132 (.ZN(net132),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_133 (.ZN(net133),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_134 (.ZN(net134),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_135 (.ZN(net135),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_136 (.ZN(net136),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_137 (.ZN(net137),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_138 (.ZN(net138),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_139 (.ZN(net139),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_140 (.ZN(net140),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_141 (.ZN(net141),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_142 (.ZN(net142),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_143 (.ZN(net143),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_144 (.ZN(net144),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_145 (.ZN(net145),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_146 (.ZN(net146),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_147 (.ZN(net147),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_148 (.ZN(net148),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_149 (.ZN(net149),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_150 (.ZN(net150),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_151 (.ZN(net151),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_152 (.ZN(net152),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_153 (.ZN(net153),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_154 (.ZN(net154),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_155 (.ZN(net155),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_156 (.ZN(net156),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_157 (.ZN(net157),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_158 (.ZN(net158),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_159 (.ZN(net159),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_160 (.ZN(net160),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_161 (.ZN(net161),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_162 (.ZN(net162),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_163 (.ZN(net163),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_164 (.ZN(net164),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_165 (.ZN(net165),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_166 (.ZN(net166),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_167 (.ZN(net167),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_168 (.ZN(net168),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_169 (.ZN(net169),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_170 (.ZN(net170),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_171 (.ZN(net171),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_172 (.ZN(net172),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_173 (.ZN(net173),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_174 (.ZN(net174),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_175 (.ZN(net175),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_176 (.ZN(net176),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_177 (.ZN(net177),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_178 (.ZN(net178),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_179 (.ZN(net179),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_180 (.ZN(net180),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_181 (.ZN(net181),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_182 (.ZN(net182),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_183 (.ZN(net183),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_184 (.ZN(net184),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_185 (.ZN(net185),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_186 (.ZN(net186),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_187 (.ZN(net187),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_188 (.ZN(net188),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_189 (.ZN(net189),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_190 (.ZN(net190),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_191 (.ZN(net191),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_192 (.ZN(net192),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_193 (.ZN(net193),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_194 (.ZN(net194),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_195 (.ZN(net195),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_196 (.ZN(net196),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_197 (.ZN(net197),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_198 (.ZN(net198),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_199 (.ZN(net199),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_200 (.ZN(net200),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_201 (.ZN(net201),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_202 (.ZN(net202),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_203 (.ZN(net203),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_204 (.ZN(net204),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_205 (.ZN(net205),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_206 (.ZN(net206),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_207 (.ZN(net207),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_208 (.ZN(net208),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_209 (.ZN(net209),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_210 (.ZN(net210),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_211 (.ZN(net211),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1 (.I(io_in[2]),
    .Z(net1),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input2 (.I(io_in[3]),
    .Z(net2),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(wb_clk_i),
    .Z(net3),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input4 (.I(wb_rst_i),
    .Z(net4),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input5 (.I(wbs_adr_i[0]),
    .Z(net5),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input6 (.I(wbs_adr_i[1]),
    .Z(net6),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input7 (.I(wbs_adr_i[2]),
    .Z(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input8 (.I(wbs_adr_i[3]),
    .Z(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input9 (.I(wbs_adr_i[4]),
    .Z(net9),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input10 (.I(wbs_adr_i[5]),
    .Z(net10),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input11 (.I(wbs_adr_i[6]),
    .Z(net11),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input12 (.I(wbs_adr_i[7]),
    .Z(net12),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input13 (.I(wbs_cyc_i),
    .Z(net13),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input14 (.I(wbs_dat_i[0]),
    .Z(net14),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input15 (.I(wbs_dat_i[10]),
    .Z(net15),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input16 (.I(wbs_dat_i[11]),
    .Z(net16),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input17 (.I(wbs_dat_i[12]),
    .Z(net17),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input18 (.I(wbs_dat_i[13]),
    .Z(net18),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input19 (.I(wbs_dat_i[14]),
    .Z(net19),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input20 (.I(wbs_dat_i[15]),
    .Z(net20),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input21 (.I(wbs_dat_i[1]),
    .Z(net21),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input22 (.I(wbs_dat_i[2]),
    .Z(net22),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input23 (.I(wbs_dat_i[3]),
    .Z(net23),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input24 (.I(wbs_dat_i[4]),
    .Z(net24),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input25 (.I(wbs_dat_i[5]),
    .Z(net25),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input26 (.I(wbs_dat_i[6]),
    .Z(net26),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input27 (.I(wbs_dat_i[7]),
    .Z(net27),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input28 (.I(wbs_dat_i[8]),
    .Z(net28),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input29 (.I(wbs_dat_i[9]),
    .Z(net29),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input30 (.I(wbs_stb_i),
    .Z(net30),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input31 (.I(wbs_we_i),
    .Z(net31),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[0]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(io_out[1]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[2]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(wbs_ack_o),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(wbs_dat_o[0]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(wbs_dat_o[10]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(wbs_dat_o[11]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(wbs_dat_o[12]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(wbs_dat_o[13]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(wbs_dat_o[14]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(wbs_dat_o[15]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(wbs_dat_o[16]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(wbs_dat_o[17]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(wbs_dat_o[18]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output46 (.I(net46),
    .Z(wbs_dat_o[19]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output47 (.I(net47),
    .Z(wbs_dat_o[1]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output48 (.I(net48),
    .Z(wbs_dat_o[20]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output49 (.I(net49),
    .Z(wbs_dat_o[21]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output50 (.I(net50),
    .Z(wbs_dat_o[22]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output51 (.I(net51),
    .Z(wbs_dat_o[23]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output52 (.I(net52),
    .Z(wbs_dat_o[24]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output53 (.I(net53),
    .Z(wbs_dat_o[25]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output54 (.I(net54),
    .Z(wbs_dat_o[26]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output55 (.I(net55),
    .Z(wbs_dat_o[27]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output56 (.I(net56),
    .Z(wbs_dat_o[28]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output57 (.I(net57),
    .Z(wbs_dat_o[29]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output58 (.I(net58),
    .Z(wbs_dat_o[2]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output59 (.I(net59),
    .Z(wbs_dat_o[30]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output60 (.I(net60),
    .Z(wbs_dat_o[31]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output61 (.I(net61),
    .Z(wbs_dat_o[3]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output62 (.I(net62),
    .Z(wbs_dat_o[4]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output63 (.I(net63),
    .Z(wbs_dat_o[5]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output64 (.I(net64),
    .Z(wbs_dat_o[6]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output65 (.I(net65),
    .Z(wbs_dat_o[7]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output66 (.I(net66),
    .Z(wbs_dat_o[8]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output67 (.I(net67),
    .Z(wbs_dat_o[9]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout68 (.I(net3),
    .Z(net68),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout69 (.I(net3),
    .Z(net69),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout70 (.I(net71),
    .Z(net70),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout71 (.I(net3),
    .Z(net71),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_project_wrapper_72 (.ZN(net72),
    .VDD(vdd),
    .VSS(vss));
 assign io_oeb[0] = net72;
 assign io_oeb[10] = net82;
 assign io_oeb[11] = net83;
 assign io_oeb[12] = net84;
 assign io_oeb[13] = net85;
 assign io_oeb[14] = net86;
 assign io_oeb[15] = net87;
 assign io_oeb[16] = net88;
 assign io_oeb[17] = net89;
 assign io_oeb[18] = net90;
 assign io_oeb[19] = net91;
 assign io_oeb[1] = net73;
 assign io_oeb[20] = net92;
 assign io_oeb[21] = net93;
 assign io_oeb[22] = net94;
 assign io_oeb[23] = net95;
 assign io_oeb[24] = net96;
 assign io_oeb[25] = net97;
 assign io_oeb[26] = net98;
 assign io_oeb[27] = net99;
 assign io_oeb[28] = net100;
 assign io_oeb[29] = net101;
 assign io_oeb[2] = net74;
 assign io_oeb[30] = net102;
 assign io_oeb[31] = net103;
 assign io_oeb[32] = net104;
 assign io_oeb[33] = net105;
 assign io_oeb[34] = net106;
 assign io_oeb[35] = net107;
 assign io_oeb[36] = net108;
 assign io_oeb[37] = net109;
 assign io_oeb[3] = net75;
 assign io_oeb[4] = net76;
 assign io_oeb[5] = net77;
 assign io_oeb[6] = net78;
 assign io_oeb[7] = net79;
 assign io_oeb[8] = net80;
 assign io_oeb[9] = net81;
 assign io_out[10] = net117;
 assign io_out[11] = net118;
 assign io_out[12] = net119;
 assign io_out[13] = net120;
 assign io_out[14] = net121;
 assign io_out[15] = net122;
 assign io_out[16] = net123;
 assign io_out[17] = net124;
 assign io_out[18] = net125;
 assign io_out[19] = net126;
 assign io_out[20] = net127;
 assign io_out[21] = net128;
 assign io_out[22] = net129;
 assign io_out[23] = net130;
 assign io_out[24] = net131;
 assign io_out[25] = net132;
 assign io_out[26] = net133;
 assign io_out[27] = net134;
 assign io_out[28] = net135;
 assign io_out[29] = net136;
 assign io_out[30] = net137;
 assign io_out[31] = net138;
 assign io_out[32] = net139;
 assign io_out[33] = net140;
 assign io_out[34] = net141;
 assign io_out[35] = net142;
 assign io_out[36] = net143;
 assign io_out[37] = net144;
 assign io_out[3] = net110;
 assign io_out[4] = net111;
 assign io_out[5] = net112;
 assign io_out[6] = net113;
 assign io_out[7] = net114;
 assign io_out[8] = net115;
 assign io_out[9] = net116;
 assign la_data_out[0] = net145;
 assign la_data_out[10] = net155;
 assign la_data_out[11] = net156;
 assign la_data_out[12] = net157;
 assign la_data_out[13] = net158;
 assign la_data_out[14] = net159;
 assign la_data_out[15] = net160;
 assign la_data_out[16] = net161;
 assign la_data_out[17] = net162;
 assign la_data_out[18] = net163;
 assign la_data_out[19] = net164;
 assign la_data_out[1] = net146;
 assign la_data_out[20] = net165;
 assign la_data_out[21] = net166;
 assign la_data_out[22] = net167;
 assign la_data_out[23] = net168;
 assign la_data_out[24] = net169;
 assign la_data_out[25] = net170;
 assign la_data_out[26] = net171;
 assign la_data_out[27] = net172;
 assign la_data_out[28] = net173;
 assign la_data_out[29] = net174;
 assign la_data_out[2] = net147;
 assign la_data_out[30] = net175;
 assign la_data_out[31] = net176;
 assign la_data_out[32] = net177;
 assign la_data_out[33] = net178;
 assign la_data_out[34] = net179;
 assign la_data_out[35] = net180;
 assign la_data_out[36] = net181;
 assign la_data_out[37] = net182;
 assign la_data_out[38] = net183;
 assign la_data_out[39] = net184;
 assign la_data_out[3] = net148;
 assign la_data_out[40] = net185;
 assign la_data_out[41] = net186;
 assign la_data_out[42] = net187;
 assign la_data_out[43] = net188;
 assign la_data_out[44] = net189;
 assign la_data_out[45] = net190;
 assign la_data_out[46] = net191;
 assign la_data_out[47] = net192;
 assign la_data_out[48] = net193;
 assign la_data_out[49] = net194;
 assign la_data_out[4] = net149;
 assign la_data_out[50] = net195;
 assign la_data_out[51] = net196;
 assign la_data_out[52] = net197;
 assign la_data_out[53] = net198;
 assign la_data_out[54] = net199;
 assign la_data_out[55] = net200;
 assign la_data_out[56] = net201;
 assign la_data_out[57] = net202;
 assign la_data_out[58] = net203;
 assign la_data_out[59] = net204;
 assign la_data_out[5] = net150;
 assign la_data_out[60] = net205;
 assign la_data_out[61] = net206;
 assign la_data_out[62] = net207;
 assign la_data_out[63] = net208;
 assign la_data_out[6] = net151;
 assign la_data_out[7] = net152;
 assign la_data_out[8] = net153;
 assign la_data_out[9] = net154;
 assign user_irq[0] = net209;
 assign user_irq[1] = net210;
 assign user_irq[2] = net211;
endmodule
