magic
tech sky130A
magscale 1 2
timestamp 1671619108
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 14 1300 59970 57712
<< metal2 >>
rect 1306 59200 1362 59800
rect 30930 59200 30986 59800
rect 59910 59200 59966 59800
rect 18 200 74 800
rect 28998 200 29054 800
rect 58622 200 58678 800
<< obsm2 >>
rect 20 59144 1250 59200
rect 1418 59144 30874 59200
rect 31042 59144 59854 59200
rect 20 856 59964 59144
rect 130 800 28942 856
rect 29110 800 58566 856
rect 58734 800 59964 856
<< metal3 >>
rect 200 30608 800 30728
rect 59200 29248 59800 29368
<< obsm3 >>
rect 800 30808 59200 57697
rect 880 30528 59200 30808
rect 800 29448 59200 30528
rect 800 29168 59120 29448
rect 800 2143 59200 29168
<< metal4 >>
rect 4208 2128 4528 57712
rect 4868 2128 5188 57712
rect 34928 2128 35248 57712
rect 35588 2128 35908 57712
<< obsm4 >>
rect 32443 26011 34848 47429
rect 35328 26011 35508 47429
rect 35988 26011 48701 47429
<< metal5 >>
rect 1056 36642 58928 36962
rect 1056 35982 58928 36302
rect 1056 6006 58928 6326
rect 1056 5346 58928 5666
<< labels >>
rlabel metal2 s 59910 59200 59966 59800 6 A_PAD
port 1 nsew signal input
rlabel metal2 s 28998 200 29054 800 6 B_PAD
port 2 nsew signal input
rlabel metal3 s 59200 29248 59800 29368 6 OUT_1
port 3 nsew signal output
rlabel metal3 s 200 30608 800 30728 6 OUT_2
port 4 nsew signal output
rlabel metal2 s 18 200 74 800 6 sel
port 5 nsew signal input
rlabel metal2 s 1306 59200 1362 59800 6 user_clock2
port 6 nsew signal input
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 7 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 7 nsew power bidirectional
rlabel metal5 s 1056 5346 58928 5666 6 vccd1
port 7 nsew power bidirectional
rlabel metal5 s 1056 35982 58928 36302 6 vccd1
port 7 nsew power bidirectional
rlabel metal4 s 4868 2128 5188 57712 6 vssd1
port 8 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 57712 6 vssd1
port 8 nsew ground bidirectional
rlabel metal5 s 1056 6006 58928 6326 6 vssd1
port 8 nsew ground bidirectional
rlabel metal5 s 1056 36642 58928 36962 6 vssd1
port 8 nsew ground bidirectional
rlabel metal2 s 30930 59200 30986 59800 6 wb_clk_i
port 9 nsew signal input
rlabel metal2 s 58622 200 58678 800 6 wb_rst_i
port 10 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3744986
string GDS_FILE /home/shahid/caravel_user_project/openlane/user_proj_asic/runs/22_12_21_15_35/results/signoff/user_proj_asic.magic.gds
string GDS_START 577154
<< end >>

