// This is the unpowered netlist.
module user_proj_asic (A_PAD,
    B_PAD,
    OUT_1,
    OUT_2,
    sel,
    user_clock2,
    wb_clk_i,
    wb_rst_i);
 input A_PAD;
 input B_PAD;
 output OUT_1;
 output OUT_2;
 input sel;
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;

 wire \MUL.PS_R1_inst1.LUT_inst1.i0 ;
 wire \MUL.PS_R1_inst1.LUT_inst1.i1 ;
 wire \MUL.PS_R1_inst1.LUT_inst1.i3 ;
 wire \MUL.PS_R1_inst1.LUT_inst1.i4 ;
 wire \MUL.PS_R1_inst1.LUT_inst10.I0 ;
 wire \MUL.PS_R1_inst1.LUT_inst10.I1 ;
 wire \MUL.PS_R1_inst1.LUT_inst11.I1 ;
 wire \MUL.PS_R1_inst1.LUT_inst12.I1 ;
 wire \MUL.PS_R1_inst1.LUT_inst13.I1 ;
 wire \MUL.PS_R1_inst1.LUT_inst14.I1 ;
 wire \MUL.PS_R1_inst1.LUT_inst15.I1 ;
 wire \MUL.PS_R1_inst1.LUT_inst2.I1 ;
 wire \MUL.PS_R1_inst1.LUT_inst3.I1 ;
 wire \MUL.PS_R1_inst1.LUT_inst4.I1 ;
 wire \MUL.PS_R1_inst1.LUT_inst5.I1 ;
 wire \MUL.PS_R1_inst1.LUT_inst6.I1 ;
 wire \MUL.PS_R1_inst1.LUT_inst7.I1 ;
 wire \MUL.PS_R1_inst1.LUT_inst8.I1 ;
 wire \MUL.PS_Rx_inst2.LUT_inst1.i3 ;
 wire \MUL.PS_Rx_inst2.LUT_inst1.i4 ;
 wire \MUL.PS_Rx_inst3.LUT_inst1.i3 ;
 wire \MUL.PS_Rx_inst3.LUT_inst1.i4 ;
 wire \MUL.PS_Rx_inst4.LUT_inst1.i3 ;
 wire \MUL.PS_Rx_inst4.LUT_inst1.i4 ;
 wire \MUL.PS_Rx_inst5.LUT_inst1.i3 ;
 wire \MUL.PS_Rx_inst5.LUT_inst1.i4 ;
 wire \MUL.PS_Rx_inst6.LUT_inst1.i3 ;
 wire \MUL.PS_Rx_inst6.LUT_inst1.i4 ;
 wire \MUL.PS_Rx_inst7.LUT_inst1.i3 ;
 wire \MUL.PS_Rx_inst7.LUT_inst1.i4 ;
 wire \MUL.PS_Rx_inst8.LUT_inst1.i3 ;
 wire \MUL.PS_Rx_inst8.LUT_inst1.i4 ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire \count2[0] ;
 wire \count2[1] ;
 wire \count2[2] ;
 wire \count2[3] ;
 wire \count2[4] ;
 wire \count2[5] ;
 wire \count[0] ;
 wire \count[1] ;
 wire \count[2] ;
 wire \count[3] ;
 wire \count[4] ;
 wire \count[5] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_0_net12;
 wire clknet_1_0__leaf_net12;
 wire clknet_1_1__leaf_net12;
 wire clknet_0_net8;
 wire clknet_1_0__leaf_net8;
 wire clknet_1_1__leaf_net8;
 wire net14;

 sky130_fd_sc_hd__clkbuf_1 _0799_ (.A(\count2[5] ),
    .X(_0090_));
 sky130_fd_sc_hd__clkbuf_1 _0800_ (.A(_0090_),
    .X(_0089_));
 sky130_fd_sc_hd__clkbuf_1 _0801_ (.A(\count2[4] ),
    .X(_0091_));
 sky130_fd_sc_hd__clkbuf_1 _0802_ (.A(_0091_),
    .X(_0088_));
 sky130_fd_sc_hd__inv_2 _0803_ (.A(\count2[2] ),
    .Y(_0092_));
 sky130_fd_sc_hd__nand2_1 _0804_ (.A(\count2[1] ),
    .B(\count2[0] ),
    .Y(_0093_));
 sky130_fd_sc_hd__and2_2 _0805_ (.A(\count2[1] ),
    .B(\count2[0] ),
    .X(_0094_));
 sky130_fd_sc_hd__and2_1 _0806_ (.A(\count[1] ),
    .B(\count[0] ),
    .X(_0095_));
 sky130_fd_sc_hd__a311oi_4 _0807_ (.A1(\count[3] ),
    .A2(\count[2] ),
    .A3(_0095_),
    .B1(\count[4] ),
    .C1(\count[5] ),
    .Y(_0096_));
 sky130_fd_sc_hd__or3_1 _0808_ (.A(\count2[5] ),
    .B(\count2[4] ),
    .C(_0096_),
    .X(_0097_));
 sky130_fd_sc_hd__a31o_1 _0809_ (.A1(\count2[3] ),
    .A2(\count2[2] ),
    .A3(_0094_),
    .B1(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__or2_1 _0810_ (.A(_0093_),
    .B(_0098_),
    .X(_0099_));
 sky130_fd_sc_hd__inv_2 _0811_ (.A(\count2[3] ),
    .Y(_0100_));
 sky130_fd_sc_hd__o21ai_1 _0812_ (.A1(_0092_),
    .A2(_0099_),
    .B1(_0100_),
    .Y(_0087_));
 sky130_fd_sc_hd__xnor2_1 _0813_ (.A(\count2[2] ),
    .B(_0099_),
    .Y(_0086_));
 sky130_fd_sc_hd__nor2_1 _0814_ (.A(\count2[1] ),
    .B(\count2[0] ),
    .Y(_0101_));
 sky130_fd_sc_hd__nor2_2 _0815_ (.A(_0094_),
    .B(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__mux2_1 _0816_ (.A0(_0102_),
    .A1(\count2[1] ),
    .S(_0098_),
    .X(_0103_));
 sky130_fd_sc_hd__clkbuf_1 _0817_ (.A(_0103_),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_4 _0818_ (.A(\count2[0] ),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_4 _0819_ (.A(_0104_),
    .X(_0105_));
 sky130_fd_sc_hd__nand2_1 _0820_ (.A(_0105_),
    .B(_0098_),
    .Y(_0106_));
 sky130_fd_sc_hd__o21ai_1 _0821_ (.A1(_0105_),
    .A2(_0097_),
    .B1(_0106_),
    .Y(_0084_));
 sky130_fd_sc_hd__buf_2 _0822_ (.A(\count[5] ),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_1 _0823_ (.A(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_1 _0824_ (.A(_0108_),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_1 _0825_ (.A(\count[4] ),
    .X(_0109_));
 sky130_fd_sc_hd__clkbuf_1 _0826_ (.A(_0109_),
    .X(_0082_));
 sky130_fd_sc_hd__inv_2 _0827_ (.A(_0095_),
    .Y(_0110_));
 sky130_fd_sc_hd__or2_1 _0828_ (.A(\count[1] ),
    .B(\count[0] ),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_4 _0829_ (.A(_0111_),
    .X(_0112_));
 sky130_fd_sc_hd__or3_2 _0830_ (.A(\count[3] ),
    .B(\count[2] ),
    .C(_0112_),
    .X(_0113_));
 sky130_fd_sc_hd__nor3_2 _0831_ (.A(_0107_),
    .B(\count[4] ),
    .C(_0113_),
    .Y(_0114_));
 sky130_fd_sc_hd__o21a_1 _0832_ (.A1(\count[4] ),
    .A2(_0113_),
    .B1(_0107_),
    .X(_0115_));
 sky130_fd_sc_hd__or3_1 _0833_ (.A(_0110_),
    .B(_0114_),
    .C(_0115_),
    .X(_0116_));
 sky130_fd_sc_hd__xnor2_4 _0834_ (.A(\count[2] ),
    .B(_0112_),
    .Y(_0117_));
 sky130_fd_sc_hd__nand2_1 _0835_ (.A(_0096_),
    .B(_0117_),
    .Y(_0118_));
 sky130_fd_sc_hd__nor2_2 _0836_ (.A(_0116_),
    .B(_0118_),
    .Y(_0119_));
 sky130_fd_sc_hd__or2_1 _0837_ (.A(\count[3] ),
    .B(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_1 _0838_ (.A(_0120_),
    .X(_0081_));
 sky130_fd_sc_hd__nor2_1 _0839_ (.A(_0107_),
    .B(\count[4] ),
    .Y(_0121_));
 sky130_fd_sc_hd__clkbuf_2 _0840_ (.A(\count[2] ),
    .X(_0122_));
 sky130_fd_sc_hd__a21oi_1 _0841_ (.A1(_0121_),
    .A2(_0095_),
    .B1(_0122_),
    .Y(_0123_));
 sky130_fd_sc_hd__nor2_1 _0842_ (.A(_0119_),
    .B(_0123_),
    .Y(_0080_));
 sky130_fd_sc_hd__a311o_1 _0843_ (.A1(\count[3] ),
    .A2(\count[2] ),
    .A3(_0095_),
    .B1(\count[4] ),
    .C1(net14),
    .X(_0124_));
 sky130_fd_sc_hd__a32o_1 _0844_ (.A1(_0121_),
    .A2(_0110_),
    .A3(_0112_),
    .B1(_0124_),
    .B2(\count[1] ),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _0845_ (.A0(_0121_),
    .A1(_0124_),
    .S(\count[0] ),
    .X(_0125_));
 sky130_fd_sc_hd__clkbuf_1 _0846_ (.A(_0125_),
    .X(_0078_));
 sky130_fd_sc_hd__clkbuf_1 _0847_ (.A(\MUL.PS_Rx_inst8.LUT_inst1.i4 ),
    .X(_0126_));
 sky130_fd_sc_hd__clkbuf_1 _0848_ (.A(_0126_),
    .X(_0075_));
 sky130_fd_sc_hd__o21ai_1 _0849_ (.A1(\count[2] ),
    .A2(_0112_),
    .B1(\count[3] ),
    .Y(_0127_));
 sky130_fd_sc_hd__a21oi_1 _0850_ (.A1(_0113_),
    .A2(_0127_),
    .B1(_0124_),
    .Y(_0128_));
 sky130_fd_sc_hd__buf_2 _0851_ (.A(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__nor3b_1 _0852_ (.A(_0107_),
    .B(\count[0] ),
    .C_N(\count[1] ),
    .Y(_0130_));
 sky130_fd_sc_hd__and2_1 _0853_ (.A(net2),
    .B(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__nand3_1 _0854_ (.A(_0122_),
    .B(_0128_),
    .C(_0130_),
    .Y(_0132_));
 sky130_fd_sc_hd__a32o_1 _0855_ (.A1(_0117_),
    .A2(_0129_),
    .A3(_0131_),
    .B1(_0132_),
    .B2(\MUL.PS_Rx_inst8.LUT_inst1.i3 ),
    .X(_0074_));
 sky130_fd_sc_hd__nor3b_1 _0856_ (.A(_0107_),
    .B(\count[1] ),
    .C_N(\count[0] ),
    .Y(_0133_));
 sky130_fd_sc_hd__and2_1 _0857_ (.A(net2),
    .B(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__nand3_1 _0858_ (.A(_0122_),
    .B(_0128_),
    .C(_0133_),
    .Y(_0135_));
 sky130_fd_sc_hd__clkbuf_4 _0859_ (.A(\MUL.PS_Rx_inst7.LUT_inst1.i4 ),
    .X(_0136_));
 sky130_fd_sc_hd__a32o_1 _0860_ (.A1(_0117_),
    .A2(_0129_),
    .A3(_0134_),
    .B1(_0135_),
    .B2(_0136_),
    .X(_0073_));
 sky130_fd_sc_hd__o21ai_1 _0861_ (.A1(\count[4] ),
    .A2(_0113_),
    .B1(_0128_),
    .Y(_0137_));
 sky130_fd_sc_hd__or3b_1 _0862_ (.A(_0112_),
    .B(_0107_),
    .C_N(\count[2] ),
    .X(_0138_));
 sky130_fd_sc_hd__nor2_1 _0863_ (.A(_0137_),
    .B(_0138_),
    .Y(_0139_));
 sky130_fd_sc_hd__mux2_1 _0864_ (.A0(\MUL.PS_Rx_inst7.LUT_inst1.i3 ),
    .A1(net2),
    .S(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_1 _0865_ (.A(_0140_),
    .X(_0072_));
 sky130_fd_sc_hd__clkbuf_4 _0866_ (.A(\MUL.PS_Rx_inst6.LUT_inst1.i4 ),
    .X(_0141_));
 sky130_fd_sc_hd__or3_1 _0867_ (.A(_0122_),
    .B(_0116_),
    .C(_0137_),
    .X(_0142_));
 sky130_fd_sc_hd__and3b_1 _0868_ (.A_N(_0107_),
    .B(\count[1] ),
    .C(\count[0] ),
    .X(_0143_));
 sky130_fd_sc_hd__xor2_4 _0869_ (.A(\count[2] ),
    .B(_0112_),
    .X(_0144_));
 sky130_fd_sc_hd__and3_1 _0870_ (.A(net2),
    .B(_0143_),
    .C(_0144_),
    .X(_0145_));
 sky130_fd_sc_hd__a22o_1 _0871_ (.A1(_0141_),
    .A2(_0142_),
    .B1(_0145_),
    .B2(_0129_),
    .X(_0071_));
 sky130_fd_sc_hd__or3b_1 _0872_ (.A(_0107_),
    .B(\count[0] ),
    .C_N(\count[1] ),
    .X(_0146_));
 sky130_fd_sc_hd__or3_1 _0873_ (.A(_0122_),
    .B(_0137_),
    .C(_0146_),
    .X(_0147_));
 sky130_fd_sc_hd__a32o_1 _0874_ (.A1(_0144_),
    .A2(_0129_),
    .A3(_0131_),
    .B1(_0147_),
    .B2(\MUL.PS_Rx_inst6.LUT_inst1.i3 ),
    .X(_0070_));
 sky130_fd_sc_hd__or3b_1 _0875_ (.A(_0107_),
    .B(\count[1] ),
    .C_N(\count[0] ),
    .X(_0148_));
 sky130_fd_sc_hd__or3_1 _0876_ (.A(\count[2] ),
    .B(_0137_),
    .C(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_4 _0877_ (.A(\MUL.PS_Rx_inst5.LUT_inst1.i4 ),
    .X(_0150_));
 sky130_fd_sc_hd__a32o_1 _0878_ (.A1(_0144_),
    .A2(_0129_),
    .A3(_0134_),
    .B1(_0149_),
    .B2(_0150_),
    .X(_0069_));
 sky130_fd_sc_hd__or4_1 _0879_ (.A(_0112_),
    .B(_0114_),
    .C(_0115_),
    .D(_0118_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _0880_ (.A0(net2),
    .A1(\MUL.PS_Rx_inst5.LUT_inst1.i3 ),
    .S(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_1 _0881_ (.A(_0152_),
    .X(_0068_));
 sky130_fd_sc_hd__clkbuf_4 _0882_ (.A(\MUL.PS_Rx_inst4.LUT_inst1.i4 ),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _0883_ (.A0(_0153_),
    .A1(net2),
    .S(_0119_),
    .X(_0154_));
 sky130_fd_sc_hd__clkbuf_1 _0884_ (.A(_0154_),
    .X(_0067_));
 sky130_fd_sc_hd__and3_1 _0885_ (.A(_0096_),
    .B(_0113_),
    .C(_0127_),
    .X(_0155_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0886_ (.A(_0155_),
    .X(_0156_));
 sky130_fd_sc_hd__buf_2 _0887_ (.A(_0156_),
    .X(_0157_));
 sky130_fd_sc_hd__nand3_1 _0888_ (.A(_0122_),
    .B(_0130_),
    .C(_0156_),
    .Y(_0158_));
 sky130_fd_sc_hd__a32o_1 _0889_ (.A1(_0117_),
    .A2(_0131_),
    .A3(_0157_),
    .B1(_0158_),
    .B2(\MUL.PS_Rx_inst4.LUT_inst1.i3 ),
    .X(_0066_));
 sky130_fd_sc_hd__nand3_1 _0890_ (.A(_0122_),
    .B(_0133_),
    .C(_0156_),
    .Y(_0159_));
 sky130_fd_sc_hd__buf_2 _0891_ (.A(\MUL.PS_Rx_inst3.LUT_inst1.i4 ),
    .X(_0160_));
 sky130_fd_sc_hd__a32o_1 _0892_ (.A1(_0117_),
    .A2(_0134_),
    .A3(_0157_),
    .B1(_0159_),
    .B2(_0160_),
    .X(_0065_));
 sky130_fd_sc_hd__and2b_1 _0893_ (.A_N(_0138_),
    .B(_0156_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _0894_ (.A0(\MUL.PS_Rx_inst3.LUT_inst1.i3 ),
    .A1(net2),
    .S(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__clkbuf_1 _0895_ (.A(_0162_),
    .X(_0064_));
 sky130_fd_sc_hd__or3b_1 _0896_ (.A(_0122_),
    .B(_0116_),
    .C_N(_0156_),
    .X(_0163_));
 sky130_fd_sc_hd__clkbuf_4 _0897_ (.A(\MUL.PS_Rx_inst2.LUT_inst1.i4 ),
    .X(_0164_));
 sky130_fd_sc_hd__a22o_1 _0898_ (.A1(_0145_),
    .A2(_0157_),
    .B1(_0163_),
    .B2(_0164_),
    .X(_0063_));
 sky130_fd_sc_hd__or3b_1 _0899_ (.A(_0122_),
    .B(_0146_),
    .C_N(_0156_),
    .X(_0165_));
 sky130_fd_sc_hd__a32o_1 _0900_ (.A1(_0144_),
    .A2(_0131_),
    .A3(_0157_),
    .B1(_0165_),
    .B2(\MUL.PS_Rx_inst2.LUT_inst1.i3 ),
    .X(_0062_));
 sky130_fd_sc_hd__or3b_1 _0901_ (.A(_0122_),
    .B(_0148_),
    .C_N(_0156_),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_4 _0902_ (.A(\MUL.PS_R1_inst1.LUT_inst1.i4 ),
    .X(_0167_));
 sky130_fd_sc_hd__a32o_1 _0903_ (.A1(_0144_),
    .A2(_0134_),
    .A3(_0157_),
    .B1(_0166_),
    .B2(_0167_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0904_ (.A0(\MUL.PS_R1_inst1.LUT_inst1.i3 ),
    .A1(net2),
    .S(_0114_),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_1 _0905_ (.A(_0168_),
    .X(_0060_));
 sky130_fd_sc_hd__buf_2 _0906_ (.A(\MUL.PS_R1_inst1.LUT_inst15.I1 ),
    .X(_0169_));
 sky130_fd_sc_hd__clkbuf_4 _0907_ (.A(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_1 _0908_ (.A(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__clkbuf_1 _0909_ (.A(_0171_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _0910_ (.A(net1),
    .B(_0130_),
    .X(_0172_));
 sky130_fd_sc_hd__buf_2 _0911_ (.A(\MUL.PS_R1_inst1.LUT_inst14.I1 ),
    .X(_0173_));
 sky130_fd_sc_hd__buf_2 _0912_ (.A(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__a32o_1 _0913_ (.A1(_0117_),
    .A2(_0129_),
    .A3(_0172_),
    .B1(_0132_),
    .B2(_0174_),
    .X(_0058_));
 sky130_fd_sc_hd__and2_1 _0914_ (.A(net1),
    .B(_0133_),
    .X(_0175_));
 sky130_fd_sc_hd__clkbuf_4 _0915_ (.A(\MUL.PS_R1_inst1.LUT_inst13.I1 ),
    .X(_0176_));
 sky130_fd_sc_hd__clkbuf_4 _0916_ (.A(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__a32o_1 _0917_ (.A1(_0117_),
    .A2(_0129_),
    .A3(_0175_),
    .B1(_0135_),
    .B2(_0177_),
    .X(_0057_));
 sky130_fd_sc_hd__buf_2 _0918_ (.A(\MUL.PS_R1_inst1.LUT_inst12.I1 ),
    .X(_0178_));
 sky130_fd_sc_hd__clkbuf_4 _0919_ (.A(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _0920_ (.A0(_0179_),
    .A1(net1),
    .S(_0139_),
    .X(_0180_));
 sky130_fd_sc_hd__clkbuf_1 _0921_ (.A(_0180_),
    .X(_0056_));
 sky130_fd_sc_hd__buf_2 _0922_ (.A(\MUL.PS_R1_inst1.LUT_inst11.I1 ),
    .X(_0181_));
 sky130_fd_sc_hd__clkbuf_4 _0923_ (.A(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__and3_1 _0924_ (.A(net1),
    .B(_0143_),
    .C(_0144_),
    .X(_0183_));
 sky130_fd_sc_hd__a22o_1 _0925_ (.A1(_0182_),
    .A2(_0142_),
    .B1(_0183_),
    .B2(_0129_),
    .X(_0055_));
 sky130_fd_sc_hd__clkbuf_4 _0926_ (.A(\MUL.PS_R1_inst1.LUT_inst10.I1 ),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_4 _0927_ (.A(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__a32o_1 _0928_ (.A1(_0144_),
    .A2(_0129_),
    .A3(_0172_),
    .B1(_0147_),
    .B2(_0185_),
    .X(_0054_));
 sky130_fd_sc_hd__clkbuf_4 _0929_ (.A(\MUL.PS_R1_inst1.LUT_inst10.I0 ),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_4 _0930_ (.A(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__a32o_1 _0931_ (.A1(_0144_),
    .A2(_0129_),
    .A3(_0175_),
    .B1(_0149_),
    .B2(_0187_),
    .X(_0053_));
 sky130_fd_sc_hd__clkbuf_4 _0932_ (.A(\MUL.PS_R1_inst1.LUT_inst8.I1 ),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_4 _0933_ (.A(_0188_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _0934_ (.A0(net1),
    .A1(_0189_),
    .S(_0151_),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_1 _0935_ (.A(_0190_),
    .X(_0052_));
 sky130_fd_sc_hd__clkbuf_4 _0936_ (.A(\MUL.PS_R1_inst1.LUT_inst7.I1 ),
    .X(_0191_));
 sky130_fd_sc_hd__clkbuf_4 _0937_ (.A(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _0938_ (.A0(_0192_),
    .A1(net1),
    .S(_0119_),
    .X(_0193_));
 sky130_fd_sc_hd__clkbuf_1 _0939_ (.A(_0193_),
    .X(_0051_));
 sky130_fd_sc_hd__clkbuf_4 _0940_ (.A(\MUL.PS_R1_inst1.LUT_inst6.I1 ),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_4 _0941_ (.A(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__a32o_1 _0942_ (.A1(_0117_),
    .A2(_0157_),
    .A3(_0172_),
    .B1(_0158_),
    .B2(_0195_),
    .X(_0050_));
 sky130_fd_sc_hd__clkbuf_4 _0943_ (.A(\MUL.PS_R1_inst1.LUT_inst5.I1 ),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_4 _0944_ (.A(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__a32o_1 _0945_ (.A1(_0117_),
    .A2(_0157_),
    .A3(_0175_),
    .B1(_0159_),
    .B2(_0197_),
    .X(_0049_));
 sky130_fd_sc_hd__clkbuf_4 _0946_ (.A(\MUL.PS_R1_inst1.LUT_inst4.I1 ),
    .X(_0198_));
 sky130_fd_sc_hd__buf_4 _0947_ (.A(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _0948_ (.A0(_0199_),
    .A1(net1),
    .S(_0161_),
    .X(_0200_));
 sky130_fd_sc_hd__clkbuf_1 _0949_ (.A(_0200_),
    .X(_0048_));
 sky130_fd_sc_hd__clkbuf_4 _0950_ (.A(\MUL.PS_R1_inst1.LUT_inst3.I1 ),
    .X(_0201_));
 sky130_fd_sc_hd__buf_4 _0951_ (.A(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__a22o_1 _0952_ (.A1(_0202_),
    .A2(_0163_),
    .B1(_0183_),
    .B2(_0157_),
    .X(_0047_));
 sky130_fd_sc_hd__clkbuf_4 _0953_ (.A(\MUL.PS_R1_inst1.LUT_inst2.I1 ),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_4 _0954_ (.A(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__a32o_1 _0955_ (.A1(_0144_),
    .A2(_0157_),
    .A3(_0172_),
    .B1(_0165_),
    .B2(_0204_),
    .X(_0046_));
 sky130_fd_sc_hd__clkbuf_4 _0956_ (.A(\MUL.PS_R1_inst1.LUT_inst1.i1 ),
    .X(_0205_));
 sky130_fd_sc_hd__a32o_1 _0957_ (.A1(_0144_),
    .A2(_0157_),
    .A3(_0175_),
    .B1(_0166_),
    .B2(_0205_),
    .X(_0045_));
 sky130_fd_sc_hd__clkbuf_4 _0958_ (.A(\MUL.PS_R1_inst1.LUT_inst1.i0 ),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _0959_ (.A0(_0206_),
    .A1(net1),
    .S(_0114_),
    .X(_0207_));
 sky130_fd_sc_hd__clkbuf_1 _0960_ (.A(_0207_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0961_ (.A0(net4),
    .A1(wb_clk_i),
    .S(net3),
    .X(_0208_));
 sky130_fd_sc_hd__clkbuf_4 _0962_ (.A(_0208_),
    .X(wb_clk_i));
 sky130_fd_sc_hd__clkbuf_4 _0963_ (.A(net5),
    .X(_0209_));
 sky130_fd_sc_hd__buf_4 _0964_ (.A(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__inv_2 _0965_ (.A(_0210_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _0966_ (.A(_0210_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _0967_ (.A(_0210_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _0968_ (.A(_0210_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0969_ (.A(_0210_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0970_ (.A(_0210_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _0971_ (.A(_0210_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _0972_ (.A(_0210_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _0973_ (.A(_0210_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _0974_ (.A(_0210_),
    .Y(_0009_));
 sky130_fd_sc_hd__buf_4 _0975_ (.A(_0209_),
    .X(_0211_));
 sky130_fd_sc_hd__inv_2 _0976_ (.A(_0211_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _0977_ (.A(_0211_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _0978_ (.A(_0211_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _0979_ (.A(_0211_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _0980_ (.A(_0211_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _0981_ (.A(_0211_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _0982_ (.A(_0211_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _0983_ (.A(_0211_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _0984_ (.A(_0211_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _0985_ (.A(_0211_),
    .Y(_0019_));
 sky130_fd_sc_hd__buf_4 _0986_ (.A(_0209_),
    .X(_0212_));
 sky130_fd_sc_hd__inv_2 _0987_ (.A(_0212_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _0988_ (.A(_0212_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _0989_ (.A(_0212_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _0990_ (.A(_0212_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _0991_ (.A(_0212_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _0992_ (.A(_0212_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _0993_ (.A(_0212_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _0994_ (.A(_0212_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _0995_ (.A(_0212_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _0996_ (.A(_0212_),
    .Y(_0029_));
 sky130_fd_sc_hd__buf_4 _0997_ (.A(_0209_),
    .X(_0213_));
 sky130_fd_sc_hd__inv_2 _0998_ (.A(_0213_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _0999_ (.A(_0213_),
    .Y(_0031_));
 sky130_fd_sc_hd__nor2_1 _1000_ (.A(_0209_),
    .B(_0098_),
    .Y(_0214_));
 sky130_fd_sc_hd__and2_1 _1001_ (.A(\MUL.PS_Rx_inst4.LUT_inst1.i3 ),
    .B(_0160_),
    .X(_0215_));
 sky130_fd_sc_hd__nor2_1 _1002_ (.A(\MUL.PS_Rx_inst4.LUT_inst1.i3 ),
    .B(_0160_),
    .Y(_0216_));
 sky130_fd_sc_hd__nor3_2 _1003_ (.A(\MUL.PS_Rx_inst4.LUT_inst1.i4 ),
    .B(_0215_),
    .C(_0216_),
    .Y(_0217_));
 sky130_fd_sc_hd__buf_2 _1004_ (.A(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__a21o_1 _1005_ (.A1(_0153_),
    .A2(_0216_),
    .B1(_0215_),
    .X(_0219_));
 sky130_fd_sc_hd__buf_2 _1006_ (.A(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__o21ai_2 _1007_ (.A1(\MUL.PS_Rx_inst4.LUT_inst1.i3 ),
    .A2(_0160_),
    .B1(\MUL.PS_Rx_inst4.LUT_inst1.i4 ),
    .Y(_0221_));
 sky130_fd_sc_hd__buf_2 _1008_ (.A(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__nand3_1 _1009_ (.A(\MUL.PS_Rx_inst4.LUT_inst1.i4 ),
    .B(\MUL.PS_Rx_inst4.LUT_inst1.i3 ),
    .C(_0160_),
    .Y(_0223_));
 sky130_fd_sc_hd__buf_2 _1010_ (.A(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__o21ai_1 _1011_ (.A1(_0203_),
    .A2(_0222_),
    .B1(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__a221o_1 _1012_ (.A1(_0203_),
    .A2(_0218_),
    .B1(_0220_),
    .B2(_0205_),
    .C1(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__clkinv_2 _1013_ (.A(\MUL.PS_Rx_inst3.LUT_inst1.i4 ),
    .Y(_0227_));
 sky130_fd_sc_hd__or2_1 _1014_ (.A(\MUL.PS_Rx_inst3.LUT_inst1.i3 ),
    .B(\MUL.PS_Rx_inst2.LUT_inst1.i4 ),
    .X(_0228_));
 sky130_fd_sc_hd__nand2_1 _1015_ (.A(\MUL.PS_Rx_inst3.LUT_inst1.i3 ),
    .B(_0164_),
    .Y(_0229_));
 sky130_fd_sc_hd__o21ai_2 _1016_ (.A1(_0227_),
    .A2(_0228_),
    .B1(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__clkbuf_4 _1017_ (.A(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__and3_1 _1018_ (.A(_0227_),
    .B(_0229_),
    .C(_0228_),
    .X(_0232_));
 sky130_fd_sc_hd__clkbuf_4 _1019_ (.A(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__o21ai_2 _1020_ (.A1(\MUL.PS_Rx_inst3.LUT_inst1.i3 ),
    .A2(_0164_),
    .B1(_0160_),
    .Y(_0234_));
 sky130_fd_sc_hd__clkbuf_4 _1021_ (.A(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__nand3_1 _1022_ (.A(_0160_),
    .B(\MUL.PS_Rx_inst3.LUT_inst1.i3 ),
    .C(_0164_),
    .Y(_0236_));
 sky130_fd_sc_hd__buf_2 _1023_ (.A(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__o21ai_1 _1024_ (.A1(_0198_),
    .A2(_0235_),
    .B1(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__a221o_1 _1025_ (.A1(\MUL.PS_R1_inst1.LUT_inst3.I1 ),
    .A2(_0231_),
    .B1(_0233_),
    .B2(_0199_),
    .C1(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__nand2_2 _1026_ (.A(\MUL.PS_Rx_inst2.LUT_inst1.i3 ),
    .B(\MUL.PS_R1_inst1.LUT_inst1.i4 ),
    .Y(_0240_));
 sky130_fd_sc_hd__or3b_2 _1027_ (.A(\MUL.PS_Rx_inst2.LUT_inst1.i3 ),
    .B(_0167_),
    .C_N(\MUL.PS_Rx_inst2.LUT_inst1.i4 ),
    .X(_0241_));
 sky130_fd_sc_hd__nand2_4 _1028_ (.A(_0240_),
    .B(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__buf_8 _1029_ (.A(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__o21ba_1 _1030_ (.A1(\MUL.PS_Rx_inst2.LUT_inst1.i3 ),
    .A2(\MUL.PS_R1_inst1.LUT_inst1.i4 ),
    .B1_N(\MUL.PS_Rx_inst2.LUT_inst1.i4 ),
    .X(_0244_));
 sky130_fd_sc_hd__and2_1 _1031_ (.A(_0240_),
    .B(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__buf_4 _1032_ (.A(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__buf_6 _1033_ (.A(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__buf_2 _1034_ (.A(_0240_),
    .X(_0248_));
 sky130_fd_sc_hd__o21ai_2 _1035_ (.A1(\MUL.PS_Rx_inst2.LUT_inst1.i3 ),
    .A2(_0167_),
    .B1(\MUL.PS_Rx_inst2.LUT_inst1.i4 ),
    .Y(_0249_));
 sky130_fd_sc_hd__buf_2 _1036_ (.A(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__a21oi_1 _1037_ (.A1(_0194_),
    .A2(_0248_),
    .B1(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__a221oi_4 _1038_ (.A1(\MUL.PS_R1_inst1.LUT_inst5.I1 ),
    .A2(_0243_),
    .B1(_0247_),
    .B2(_0194_),
    .C1(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__a21oi_1 _1039_ (.A1(_0196_),
    .A2(_0248_),
    .B1(_0250_),
    .Y(_0253_));
 sky130_fd_sc_hd__a221oi_4 _1040_ (.A1(_0198_),
    .A2(_0243_),
    .B1(_0247_),
    .B2(_0196_),
    .C1(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__xnor2_1 _1041_ (.A(_0252_),
    .B(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__xnor2_1 _1042_ (.A(_0239_),
    .B(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__o21ai_1 _1043_ (.A1(_0201_),
    .A2(_0235_),
    .B1(_0237_),
    .Y(_0257_));
 sky130_fd_sc_hd__a221o_1 _1044_ (.A1(\MUL.PS_R1_inst1.LUT_inst2.I1 ),
    .A2(_0231_),
    .B1(_0233_),
    .B2(_0202_),
    .C1(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__a21oi_1 _1045_ (.A1(_0198_),
    .A2(_0248_),
    .B1(_0250_),
    .Y(_0259_));
 sky130_fd_sc_hd__a221oi_4 _1046_ (.A1(_0201_),
    .A2(_0243_),
    .B1(_0247_),
    .B2(_0199_),
    .C1(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__xnor2_1 _1047_ (.A(_0254_),
    .B(_0260_),
    .Y(_0261_));
 sky130_fd_sc_hd__xnor2_2 _1048_ (.A(_0258_),
    .B(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__xor2_1 _1049_ (.A(_0256_),
    .B(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__xnor2_1 _1050_ (.A(_0226_),
    .B(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__o21ai_1 _1051_ (.A1(_0202_),
    .A2(_0222_),
    .B1(_0224_),
    .Y(_0265_));
 sky130_fd_sc_hd__a221o_1 _1052_ (.A1(_0202_),
    .A2(_0218_),
    .B1(_0220_),
    .B2(_0203_),
    .C1(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__o21ai_1 _1053_ (.A1(_0196_),
    .A2(_0235_),
    .B1(_0237_),
    .Y(_0267_));
 sky130_fd_sc_hd__a221o_1 _1054_ (.A1(\MUL.PS_R1_inst1.LUT_inst4.I1 ),
    .A2(_0231_),
    .B1(_0233_),
    .B2(_0196_),
    .C1(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__a21oi_1 _1055_ (.A1(_0191_),
    .A2(_0248_),
    .B1(_0250_),
    .Y(_0269_));
 sky130_fd_sc_hd__a221oi_4 _1056_ (.A1(\MUL.PS_R1_inst1.LUT_inst6.I1 ),
    .A2(_0243_),
    .B1(_0247_),
    .B2(_0191_),
    .C1(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__xnor2_1 _1057_ (.A(_0270_),
    .B(_0252_),
    .Y(_0271_));
 sky130_fd_sc_hd__xnor2_1 _1058_ (.A(_0268_),
    .B(_0271_),
    .Y(_0272_));
 sky130_fd_sc_hd__xnor2_1 _1059_ (.A(_0272_),
    .B(_0256_),
    .Y(_0273_));
 sky130_fd_sc_hd__xnor2_2 _1060_ (.A(_0266_),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__and2_1 _1061_ (.A(\MUL.PS_Rx_inst5.LUT_inst1.i3 ),
    .B(_0153_),
    .X(_0275_));
 sky130_fd_sc_hd__nor2_1 _1062_ (.A(\MUL.PS_Rx_inst5.LUT_inst1.i3 ),
    .B(_0153_),
    .Y(_0276_));
 sky130_fd_sc_hd__nor3_2 _1063_ (.A(\MUL.PS_Rx_inst5.LUT_inst1.i4 ),
    .B(_0275_),
    .C(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__buf_2 _1064_ (.A(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__inv_2 _1065_ (.A(_0153_),
    .Y(_0279_));
 sky130_fd_sc_hd__a21o_1 _1066_ (.A1(_0150_),
    .A2(\MUL.PS_Rx_inst5.LUT_inst1.i3 ),
    .B1(\MUL.PS_R1_inst1.LUT_inst1.i0 ),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _1067_ (.A0(_0279_),
    .A1(_0275_),
    .S(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__a21oi_1 _1068_ (.A1(\MUL.PS_R1_inst1.LUT_inst1.i1 ),
    .A2(_0278_),
    .B1(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__xnor2_1 _1069_ (.A(_0150_),
    .B(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__xnor2_1 _1070_ (.A(_0274_),
    .B(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__mux2_1 _1071_ (.A0(_0264_),
    .A1(_0284_),
    .S(_0105_),
    .X(_0285_));
 sky130_fd_sc_hd__a21o_1 _1072_ (.A1(\MUL.PS_Rx_inst5.LUT_inst1.i4 ),
    .A2(_0276_),
    .B1(_0275_),
    .X(_0286_));
 sky130_fd_sc_hd__buf_2 _1073_ (.A(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__o21ai_2 _1074_ (.A1(\MUL.PS_Rx_inst5.LUT_inst1.i3 ),
    .A2(_0153_),
    .B1(\MUL.PS_Rx_inst5.LUT_inst1.i4 ),
    .Y(_0288_));
 sky130_fd_sc_hd__buf_2 _1075_ (.A(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__nand3_2 _1076_ (.A(\MUL.PS_Rx_inst5.LUT_inst1.i4 ),
    .B(\MUL.PS_Rx_inst5.LUT_inst1.i3 ),
    .C(_0153_),
    .Y(_0290_));
 sky130_fd_sc_hd__buf_2 _1077_ (.A(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__o21ai_1 _1078_ (.A1(_0201_),
    .A2(_0289_),
    .B1(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__a221o_1 _1079_ (.A1(_0203_),
    .A2(_0287_),
    .B1(_0278_),
    .B2(_0202_),
    .C1(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__o21ai_1 _1080_ (.A1(_0196_),
    .A2(_0222_),
    .B1(_0224_),
    .Y(_0294_));
 sky130_fd_sc_hd__a221o_1 _1081_ (.A1(_0196_),
    .A2(_0218_),
    .B1(_0220_),
    .B2(\MUL.PS_R1_inst1.LUT_inst4.I1 ),
    .C1(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__a21oi_1 _1082_ (.A1(_0186_),
    .A2(_0248_),
    .B1(_0250_),
    .Y(_0296_));
 sky130_fd_sc_hd__a221oi_4 _1083_ (.A1(\MUL.PS_R1_inst1.LUT_inst8.I1 ),
    .A2(_0243_),
    .B1(_0247_),
    .B2(_0186_),
    .C1(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__o21ai_1 _1084_ (.A1(\MUL.PS_R1_inst1.LUT_inst7.I1 ),
    .A2(_0235_),
    .B1(_0237_),
    .Y(_0298_));
 sky130_fd_sc_hd__a221o_1 _1085_ (.A1(\MUL.PS_R1_inst1.LUT_inst6.I1 ),
    .A2(_0231_),
    .B1(_0233_),
    .B2(\MUL.PS_R1_inst1.LUT_inst7.I1 ),
    .C1(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__a21oi_1 _1086_ (.A1(\MUL.PS_R1_inst1.LUT_inst8.I1 ),
    .A2(_0248_),
    .B1(_0250_),
    .Y(_0300_));
 sky130_fd_sc_hd__a221oi_4 _1087_ (.A1(\MUL.PS_R1_inst1.LUT_inst7.I1 ),
    .A2(_0243_),
    .B1(_0247_),
    .B2(_0188_),
    .C1(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__xor2_1 _1088_ (.A(_0299_),
    .B(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__xnor2_1 _1089_ (.A(_0297_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__o21ai_1 _1090_ (.A1(\MUL.PS_R1_inst1.LUT_inst6.I1 ),
    .A2(_0235_),
    .B1(_0237_),
    .Y(_0304_));
 sky130_fd_sc_hd__a221o_1 _1091_ (.A1(\MUL.PS_R1_inst1.LUT_inst5.I1 ),
    .A2(_0231_),
    .B1(_0233_),
    .B2(_0194_),
    .C1(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__xor2_1 _1092_ (.A(_0301_),
    .B(_0270_),
    .X(_0306_));
 sky130_fd_sc_hd__xnor2_1 _1093_ (.A(_0305_),
    .B(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__xnor2_1 _1094_ (.A(_0303_),
    .B(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__xnor2_1 _1095_ (.A(_0295_),
    .B(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__o21ai_1 _1096_ (.A1(_0198_),
    .A2(_0222_),
    .B1(_0224_),
    .Y(_0310_));
 sky130_fd_sc_hd__a221o_1 _1097_ (.A1(_0198_),
    .A2(_0218_),
    .B1(_0220_),
    .B2(\MUL.PS_R1_inst1.LUT_inst3.I1 ),
    .C1(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__xnor2_1 _1098_ (.A(_0307_),
    .B(_0272_),
    .Y(_0312_));
 sky130_fd_sc_hd__xnor2_1 _1099_ (.A(_0311_),
    .B(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__xor2_1 _1100_ (.A(_0309_),
    .B(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__xnor2_2 _1101_ (.A(_0293_),
    .B(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__and2_1 _1102_ (.A(\MUL.PS_Rx_inst6.LUT_inst1.i3 ),
    .B(\MUL.PS_Rx_inst5.LUT_inst1.i4 ),
    .X(_0316_));
 sky130_fd_sc_hd__nor2_1 _1103_ (.A(\MUL.PS_Rx_inst6.LUT_inst1.i3 ),
    .B(_0150_),
    .Y(_0317_));
 sky130_fd_sc_hd__nor2_1 _1104_ (.A(\MUL.PS_Rx_inst6.LUT_inst1.i4 ),
    .B(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__and2b_1 _1105_ (.A_N(_0316_),
    .B(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__buf_2 _1106_ (.A(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__inv_2 _1107_ (.A(_0150_),
    .Y(_0321_));
 sky130_fd_sc_hd__a21o_1 _1108_ (.A1(_0141_),
    .A2(\MUL.PS_Rx_inst6.LUT_inst1.i3 ),
    .B1(_0206_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _1109_ (.A0(_0321_),
    .A1(_0316_),
    .S(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__a21oi_1 _1110_ (.A1(_0205_),
    .A2(_0320_),
    .B1(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__xnor2_1 _1111_ (.A(_0141_),
    .B(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__xnor2_1 _1112_ (.A(_0315_),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__o21ai_1 _1113_ (.A1(_0204_),
    .A2(_0289_),
    .B1(_0291_),
    .Y(_0327_));
 sky130_fd_sc_hd__a221o_1 _1114_ (.A1(_0205_),
    .A2(_0287_),
    .B1(_0278_),
    .B2(_0204_),
    .C1(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__xor2_1 _1115_ (.A(_0313_),
    .B(_0274_),
    .X(_0329_));
 sky130_fd_sc_hd__xnor2_1 _1116_ (.A(_0328_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__nor2_1 _1117_ (.A(_0105_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__inv_2 _1118_ (.A(\count2[1] ),
    .Y(_0332_));
 sky130_fd_sc_hd__a211o_1 _1119_ (.A1(_0105_),
    .A2(_0326_),
    .B1(_0331_),
    .C1(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__o21ai_1 _1120_ (.A1(\count2[1] ),
    .A2(_0285_),
    .B1(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__o21ai_1 _1121_ (.A1(_0188_),
    .A2(_0235_),
    .B1(_0237_),
    .Y(_0335_));
 sky130_fd_sc_hd__a221o_1 _1122_ (.A1(_0191_),
    .A2(_0231_),
    .B1(_0233_),
    .B2(_0188_),
    .C1(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__a21oi_1 _1123_ (.A1(\MUL.PS_R1_inst1.LUT_inst10.I1 ),
    .A2(_0240_),
    .B1(_0250_),
    .Y(_0337_));
 sky130_fd_sc_hd__a221oi_4 _1124_ (.A1(\MUL.PS_R1_inst1.LUT_inst10.I0 ),
    .A2(_0243_),
    .B1(_0246_),
    .B2(_0184_),
    .C1(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__xnor2_1 _1125_ (.A(_0297_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__xnor2_2 _1126_ (.A(_0336_),
    .B(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__o21ai_1 _1127_ (.A1(_0191_),
    .A2(_0221_),
    .B1(_0223_),
    .Y(_0341_));
 sky130_fd_sc_hd__a221o_1 _1128_ (.A1(_0191_),
    .A2(_0217_),
    .B1(_0219_),
    .B2(_0194_),
    .C1(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__o21ai_1 _1129_ (.A1(\MUL.PS_R1_inst1.LUT_inst10.I0 ),
    .A2(_0235_),
    .B1(_0237_),
    .Y(_0343_));
 sky130_fd_sc_hd__a221o_1 _1130_ (.A1(_0188_),
    .A2(_0231_),
    .B1(_0233_),
    .B2(_0186_),
    .C1(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__a21oi_1 _1131_ (.A1(\MUL.PS_R1_inst1.LUT_inst11.I1 ),
    .A2(_0240_),
    .B1(_0249_),
    .Y(_0345_));
 sky130_fd_sc_hd__a221oi_4 _1132_ (.A1(\MUL.PS_R1_inst1.LUT_inst10.I1 ),
    .A2(_0242_),
    .B1(_0246_),
    .B2(\MUL.PS_R1_inst1.LUT_inst11.I1 ),
    .C1(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__xor2_1 _1133_ (.A(_0338_),
    .B(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__xnor2_2 _1134_ (.A(_0344_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__xnor2_1 _1135_ (.A(_0342_),
    .B(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__xnor2_2 _1136_ (.A(_0340_),
    .B(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__a21oi_1 _1137_ (.A1(_0196_),
    .A2(_0291_),
    .B1(_0289_),
    .Y(_0351_));
 sky130_fd_sc_hd__a221o_1 _1138_ (.A1(\MUL.PS_R1_inst1.LUT_inst4.I1 ),
    .A2(_0287_),
    .B1(_0278_),
    .B2(_0196_),
    .C1(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__o21ai_1 _1139_ (.A1(_0194_),
    .A2(_0222_),
    .B1(_0224_),
    .Y(_0353_));
 sky130_fd_sc_hd__a221o_1 _1140_ (.A1(_0194_),
    .A2(_0218_),
    .B1(_0220_),
    .B2(_0196_),
    .C1(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__xor2_1 _1141_ (.A(_0340_),
    .B(_0303_),
    .X(_0355_));
 sky130_fd_sc_hd__xnor2_1 _1142_ (.A(_0354_),
    .B(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__xnor2_1 _1143_ (.A(_0352_),
    .B(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__xnor2_2 _1144_ (.A(_0350_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__o21ai_1 _1145_ (.A1(_0194_),
    .A2(_0288_),
    .B1(_0291_),
    .Y(_0359_));
 sky130_fd_sc_hd__a221o_1 _1146_ (.A1(\MUL.PS_R1_inst1.LUT_inst5.I1 ),
    .A2(_0286_),
    .B1(_0277_),
    .B2(_0194_),
    .C1(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__o21ai_1 _1147_ (.A1(\MUL.PS_R1_inst1.LUT_inst8.I1 ),
    .A2(_0221_),
    .B1(_0223_),
    .Y(_0361_));
 sky130_fd_sc_hd__a221o_1 _1148_ (.A1(_0188_),
    .A2(_0217_),
    .B1(_0219_),
    .B2(_0191_),
    .C1(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__o21ai_1 _1149_ (.A1(\MUL.PS_R1_inst1.LUT_inst10.I1 ),
    .A2(_0234_),
    .B1(_0236_),
    .Y(_0363_));
 sky130_fd_sc_hd__a221o_1 _1150_ (.A1(\MUL.PS_R1_inst1.LUT_inst10.I0 ),
    .A2(_0230_),
    .B1(_0232_),
    .B2(_0184_),
    .C1(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__a21oi_1 _1151_ (.A1(\MUL.PS_R1_inst1.LUT_inst12.I1 ),
    .A2(_0240_),
    .B1(_0249_),
    .Y(_0365_));
 sky130_fd_sc_hd__a221oi_4 _1152_ (.A1(\MUL.PS_R1_inst1.LUT_inst11.I1 ),
    .A2(_0242_),
    .B1(_0246_),
    .B2(\MUL.PS_R1_inst1.LUT_inst12.I1 ),
    .C1(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__xor2_1 _1153_ (.A(_0346_),
    .B(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__xnor2_1 _1154_ (.A(_0364_),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__xnor2_1 _1155_ (.A(_0362_),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__xnor2_2 _1156_ (.A(_0348_),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__xor2_1 _1157_ (.A(_0360_),
    .B(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__xnor2_1 _1158_ (.A(_0350_),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__a21o_1 _1159_ (.A1(\MUL.PS_Rx_inst6.LUT_inst1.i4 ),
    .A2(_0317_),
    .B1(_0316_),
    .X(_0373_));
 sky130_fd_sc_hd__buf_2 _1160_ (.A(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__nand3_2 _1161_ (.A(\MUL.PS_Rx_inst6.LUT_inst1.i4 ),
    .B(\MUL.PS_Rx_inst6.LUT_inst1.i3 ),
    .C(_0150_),
    .Y(_0375_));
 sky130_fd_sc_hd__buf_2 _1162_ (.A(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__o21ai_2 _1163_ (.A1(\MUL.PS_Rx_inst6.LUT_inst1.i3 ),
    .A2(_0150_),
    .B1(\MUL.PS_Rx_inst6.LUT_inst1.i4 ),
    .Y(_0377_));
 sky130_fd_sc_hd__buf_2 _1164_ (.A(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__a21oi_1 _1165_ (.A1(_0198_),
    .A2(_0376_),
    .B1(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__a221o_1 _1166_ (.A1(_0198_),
    .A2(_0320_),
    .B1(_0374_),
    .B2(\MUL.PS_R1_inst1.LUT_inst3.I1 ),
    .C1(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__xnor2_1 _1167_ (.A(_0372_),
    .B(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__xnor2_2 _1168_ (.A(_0358_),
    .B(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__a21oi_1 _1169_ (.A1(_0197_),
    .A2(_0376_),
    .B1(_0378_),
    .Y(_0383_));
 sky130_fd_sc_hd__a221o_1 _1170_ (.A1(_0197_),
    .A2(_0320_),
    .B1(_0374_),
    .B2(_0198_),
    .C1(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__o21ai_1 _1171_ (.A1(_0186_),
    .A2(_0222_),
    .B1(_0224_),
    .Y(_0385_));
 sky130_fd_sc_hd__a221o_1 _1172_ (.A1(_0186_),
    .A2(_0217_),
    .B1(_0220_),
    .B2(_0188_),
    .C1(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__o21ai_1 _1173_ (.A1(_0181_),
    .A2(_0234_),
    .B1(_0236_),
    .Y(_0387_));
 sky130_fd_sc_hd__a221o_1 _1174_ (.A1(_0184_),
    .A2(_0230_),
    .B1(_0232_),
    .B2(_0181_),
    .C1(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__a21oi_1 _1175_ (.A1(\MUL.PS_R1_inst1.LUT_inst13.I1 ),
    .A2(_0240_),
    .B1(_0249_),
    .Y(_0389_));
 sky130_fd_sc_hd__a221oi_4 _1176_ (.A1(\MUL.PS_R1_inst1.LUT_inst12.I1 ),
    .A2(_0242_),
    .B1(_0246_),
    .B2(_0176_),
    .C1(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__xor2_1 _1177_ (.A(_0366_),
    .B(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__xnor2_1 _1178_ (.A(_0388_),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__xnor2_1 _1179_ (.A(_0368_),
    .B(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__xnor2_2 _1180_ (.A(_0386_),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__a21oi_1 _1181_ (.A1(_0191_),
    .A2(_0290_),
    .B1(_0288_),
    .Y(_0395_));
 sky130_fd_sc_hd__a221o_1 _1182_ (.A1(_0194_),
    .A2(_0286_),
    .B1(_0277_),
    .B2(_0191_),
    .C1(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__xor2_1 _1183_ (.A(_0370_),
    .B(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__xnor2_2 _1184_ (.A(_0394_),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__xnor2_1 _1185_ (.A(_0372_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__xnor2_1 _1186_ (.A(_0384_),
    .B(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__o21ai_2 _1187_ (.A1(\MUL.PS_Rx_inst7.LUT_inst1.i3 ),
    .A2(_0141_),
    .B1(\MUL.PS_Rx_inst7.LUT_inst1.i4 ),
    .Y(_0401_));
 sky130_fd_sc_hd__clkbuf_4 _1188_ (.A(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__and2_1 _1189_ (.A(\MUL.PS_Rx_inst7.LUT_inst1.i3 ),
    .B(\MUL.PS_Rx_inst6.LUT_inst1.i4 ),
    .X(_0403_));
 sky130_fd_sc_hd__nor2_1 _1190_ (.A(\MUL.PS_Rx_inst7.LUT_inst1.i3 ),
    .B(_0141_),
    .Y(_0404_));
 sky130_fd_sc_hd__nor3_4 _1191_ (.A(\MUL.PS_Rx_inst7.LUT_inst1.i4 ),
    .B(_0403_),
    .C(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__a21o_2 _1192_ (.A1(\MUL.PS_Rx_inst7.LUT_inst1.i4 ),
    .A2(_0404_),
    .B1(_0403_),
    .X(_0406_));
 sky130_fd_sc_hd__a22oi_1 _1193_ (.A1(_0201_),
    .A2(_0405_),
    .B1(_0406_),
    .B2(\MUL.PS_R1_inst1.LUT_inst2.I1 ),
    .Y(_0407_));
 sky130_fd_sc_hd__nand3_2 _1194_ (.A(\MUL.PS_Rx_inst7.LUT_inst1.i4 ),
    .B(\MUL.PS_Rx_inst7.LUT_inst1.i3 ),
    .C(_0141_),
    .Y(_0408_));
 sky130_fd_sc_hd__buf_2 _1195_ (.A(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__o211a_1 _1196_ (.A1(_0201_),
    .A2(_0402_),
    .B1(_0407_),
    .C1(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__xnor2_1 _1197_ (.A(_0400_),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__xnor2_2 _1198_ (.A(_0382_),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__and2_1 _1199_ (.A(\MUL.PS_Rx_inst8.LUT_inst1.i3 ),
    .B(\MUL.PS_Rx_inst7.LUT_inst1.i4 ),
    .X(_0413_));
 sky130_fd_sc_hd__nor2_1 _1200_ (.A(\MUL.PS_Rx_inst8.LUT_inst1.i3 ),
    .B(_0136_),
    .Y(_0414_));
 sky130_fd_sc_hd__nor3_2 _1201_ (.A(\MUL.PS_Rx_inst8.LUT_inst1.i4 ),
    .B(_0413_),
    .C(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__buf_2 _1202_ (.A(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__inv_2 _1203_ (.A(_0136_),
    .Y(_0417_));
 sky130_fd_sc_hd__a21o_1 _1204_ (.A1(\MUL.PS_Rx_inst8.LUT_inst1.i4 ),
    .A2(\MUL.PS_Rx_inst8.LUT_inst1.i3 ),
    .B1(_0206_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _1205_ (.A0(_0417_),
    .A1(_0413_),
    .S(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__a21o_1 _1206_ (.A1(_0205_),
    .A2(_0416_),
    .B1(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__xor2_1 _1207_ (.A(\MUL.PS_Rx_inst8.LUT_inst1.i4 ),
    .B(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__xor2_1 _1208_ (.A(_0412_),
    .B(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_4 _1209_ (.A(_0405_),
    .X(_0423_));
 sky130_fd_sc_hd__buf_2 _1210_ (.A(_0406_),
    .X(_0424_));
 sky130_fd_sc_hd__o21ai_1 _1211_ (.A1(_0203_),
    .A2(_0402_),
    .B1(_0409_),
    .Y(_0425_));
 sky130_fd_sc_hd__a221o_1 _1212_ (.A1(_0203_),
    .A2(_0423_),
    .B1(_0424_),
    .B2(\MUL.PS_R1_inst1.LUT_inst1.i1 ),
    .C1(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__o21ai_1 _1213_ (.A1(_0201_),
    .A2(_0378_),
    .B1(_0376_),
    .Y(_0427_));
 sky130_fd_sc_hd__a221o_1 _1214_ (.A1(_0201_),
    .A2(_0320_),
    .B1(_0374_),
    .B2(\MUL.PS_R1_inst1.LUT_inst2.I1 ),
    .C1(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__a21oi_1 _1215_ (.A1(_0198_),
    .A2(_0291_),
    .B1(_0289_),
    .Y(_0429_));
 sky130_fd_sc_hd__a221o_1 _1216_ (.A1(_0201_),
    .A2(_0287_),
    .B1(_0278_),
    .B2(_0199_),
    .C1(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__xnor2_1 _1217_ (.A(_0356_),
    .B(_0309_),
    .Y(_0431_));
 sky130_fd_sc_hd__xnor2_1 _1218_ (.A(_0430_),
    .B(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__xor2_1 _1219_ (.A(_0428_),
    .B(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__xnor2_2 _1220_ (.A(_0358_),
    .B(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__xnor2_1 _1221_ (.A(_0426_),
    .B(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__xnor2_1 _1222_ (.A(_0382_),
    .B(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__xnor2_1 _1223_ (.A(_0432_),
    .B(_0315_),
    .Y(_0437_));
 sky130_fd_sc_hd__a21oi_1 _1224_ (.A1(_0203_),
    .A2(_0376_),
    .B1(_0378_),
    .Y(_0438_));
 sky130_fd_sc_hd__a221o_1 _1225_ (.A1(_0204_),
    .A2(_0320_),
    .B1(_0374_),
    .B2(_0205_),
    .C1(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__xnor2_1 _1226_ (.A(_0437_),
    .B(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__nor2_1 _1227_ (.A(\count2[1] ),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__a211o_1 _1228_ (.A1(\count2[1] ),
    .A2(_0436_),
    .B1(_0441_),
    .C1(_0105_),
    .X(_0442_));
 sky130_fd_sc_hd__inv_2 _1229_ (.A(_0141_),
    .Y(_0443_));
 sky130_fd_sc_hd__a21o_1 _1230_ (.A1(_0136_),
    .A2(\MUL.PS_Rx_inst7.LUT_inst1.i3 ),
    .B1(\MUL.PS_R1_inst1.LUT_inst1.i0 ),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _1231_ (.A0(_0443_),
    .A1(_0403_),
    .S(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__a21o_1 _1232_ (.A1(\MUL.PS_R1_inst1.LUT_inst1.i1 ),
    .A2(_0423_),
    .B1(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__xnor2_1 _1233_ (.A(_0136_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__xnor2_1 _1234_ (.A(_0434_),
    .B(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__and2_1 _1235_ (.A(_0332_),
    .B(\count2[0] ),
    .X(_0449_));
 sky130_fd_sc_hd__a21oi_1 _1236_ (.A1(_0448_),
    .A2(_0449_),
    .B1(_0092_),
    .Y(_0450_));
 sky130_fd_sc_hd__o211ai_1 _1237_ (.A1(_0093_),
    .A2(_0422_),
    .B1(_0442_),
    .C1(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__o211a_1 _1238_ (.A1(\count2[2] ),
    .A2(_0334_),
    .B1(_0451_),
    .C1(\count2[3] ),
    .X(_0452_));
 sky130_fd_sc_hd__a21o_1 _1239_ (.A1(_0153_),
    .A2(\MUL.PS_Rx_inst4.LUT_inst1.i3 ),
    .B1(_0206_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _1240_ (.A0(_0227_),
    .A1(_0215_),
    .S(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__a21oi_1 _1241_ (.A1(\MUL.PS_R1_inst1.LUT_inst1.i1 ),
    .A2(_0218_),
    .B1(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__xnor2_1 _1242_ (.A(_0279_),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__xnor2_1 _1243_ (.A(_0262_),
    .B(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__o21ai_1 _1244_ (.A1(_0203_),
    .A2(_0235_),
    .B1(_0237_),
    .Y(_0458_));
 sky130_fd_sc_hd__a221o_1 _1245_ (.A1(_0205_),
    .A2(_0231_),
    .B1(_0233_),
    .B2(_0204_),
    .C1(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__a21oi_1 _1246_ (.A1(_0202_),
    .A2(_0248_),
    .B1(_0250_),
    .Y(_0460_));
 sky130_fd_sc_hd__a221oi_4 _1247_ (.A1(_0203_),
    .A2(_0243_),
    .B1(_0247_),
    .B2(_0202_),
    .C1(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__xnor2_1 _1248_ (.A(_0260_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__xnor2_1 _1249_ (.A(_0459_),
    .B(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__nor2_1 _1250_ (.A(_0332_),
    .B(_0104_),
    .Y(_0464_));
 sky130_fd_sc_hd__a21o_1 _1251_ (.A1(_0160_),
    .A2(\MUL.PS_Rx_inst3.LUT_inst1.i3 ),
    .B1(_0206_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _1252_ (.A0(_0164_),
    .A1(_0229_),
    .S(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__a21bo_1 _1253_ (.A1(_0205_),
    .A2(_0233_),
    .B1_N(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__xnor2_1 _1254_ (.A(_0227_),
    .B(_0461_),
    .Y(_0468_));
 sky130_fd_sc_hd__xnor2_1 _1255_ (.A(_0467_),
    .B(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__a21oi_1 _1256_ (.A1(_0204_),
    .A2(_0248_),
    .B1(_0250_),
    .Y(_0470_));
 sky130_fd_sc_hd__a221o_1 _1257_ (.A1(_0205_),
    .A2(_0243_),
    .B1(_0247_),
    .B2(_0204_),
    .C1(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__a221o_1 _1258_ (.A1(_0449_),
    .A2(_0469_),
    .B1(_0471_),
    .B2(_0101_),
    .C1(_0092_),
    .X(_0472_));
 sky130_fd_sc_hd__a221o_1 _1259_ (.A1(_0094_),
    .A2(_0457_),
    .B1(_0463_),
    .B2(_0464_),
    .C1(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__inv_2 _1260_ (.A(\MUL.PS_R1_inst1.LUT_inst1.i1 ),
    .Y(_0474_));
 sky130_fd_sc_hd__o21ai_1 _1261_ (.A1(_0474_),
    .A2(_0206_),
    .B1(\MUL.PS_R1_inst1.LUT_inst1.i3 ),
    .Y(_0475_));
 sky130_fd_sc_hd__and2_1 _1262_ (.A(_0167_),
    .B(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__nor2_1 _1263_ (.A(_0164_),
    .B(_0206_),
    .Y(_0477_));
 sky130_fd_sc_hd__o211a_2 _1264_ (.A1(_0474_),
    .A2(\MUL.PS_R1_inst1.LUT_inst1.i0 ),
    .B1(_0167_),
    .C1(\MUL.PS_R1_inst1.LUT_inst1.i3 ),
    .X(_0478_));
 sky130_fd_sc_hd__inv_2 _1265_ (.A(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__o21ai_1 _1266_ (.A1(_0167_),
    .A2(_0477_),
    .B1(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__nand2_1 _1267_ (.A(\MUL.PS_R1_inst1.LUT_inst1.i1 ),
    .B(_0247_),
    .Y(_0481_));
 sky130_fd_sc_hd__o221a_1 _1268_ (.A1(_0206_),
    .A2(_0241_),
    .B1(_0477_),
    .B2(_0248_),
    .C1(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _1269_ (.A0(_0476_),
    .A1(_0480_),
    .S(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__xnor2_1 _1270_ (.A(_0164_),
    .B(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__nor2_1 _1271_ (.A(_0167_),
    .B(_0475_),
    .Y(_0485_));
 sky130_fd_sc_hd__or2_1 _1272_ (.A(_0476_),
    .B(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__a221o_1 _1273_ (.A1(_0206_),
    .A2(_0101_),
    .B1(_0464_),
    .B2(_0476_),
    .C1(\count2[2] ),
    .X(_0487_));
 sky130_fd_sc_hd__a21o_1 _1274_ (.A1(_0449_),
    .A2(_0486_),
    .B1(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__a21o_1 _1275_ (.A1(_0094_),
    .A2(_0484_),
    .B1(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__a311o_1 _1276_ (.A1(_0100_),
    .A2(_0473_),
    .A3(_0489_),
    .B1(net5),
    .C1(_0098_),
    .X(_0490_));
 sky130_fd_sc_hd__o22a_1 _1277_ (.A1(net6),
    .A2(_0214_),
    .B1(_0452_),
    .B2(_0490_),
    .X(_0076_));
 sky130_fd_sc_hd__nand2_1 _1278_ (.A(_0092_),
    .B(_0101_),
    .Y(_0491_));
 sky130_fd_sc_hd__or2_1 _1279_ (.A(\count2[1] ),
    .B(\count2[0] ),
    .X(_0492_));
 sky130_fd_sc_hd__nand2_1 _1280_ (.A(\count2[2] ),
    .B(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__nand2_1 _1281_ (.A(_0491_),
    .B(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__a21o_1 _1282_ (.A1(\MUL.PS_Rx_inst8.LUT_inst1.i4 ),
    .A2(_0414_),
    .B1(_0413_),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_2 _1283_ (.A(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__o21ai_2 _1284_ (.A1(\MUL.PS_Rx_inst8.LUT_inst1.i3 ),
    .A2(_0136_),
    .B1(\MUL.PS_Rx_inst8.LUT_inst1.i4 ),
    .Y(_0497_));
 sky130_fd_sc_hd__clkbuf_2 _1285_ (.A(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__nand2_1 _1286_ (.A(\MUL.PS_Rx_inst8.LUT_inst1.i4 ),
    .B(_0413_),
    .Y(_0499_));
 sky130_fd_sc_hd__o21ai_1 _1287_ (.A1(_0202_),
    .A2(_0498_),
    .B1(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__a221o_1 _1288_ (.A1(_0202_),
    .A2(_0416_),
    .B1(_0496_),
    .B2(_0204_),
    .C1(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__a21oi_1 _1289_ (.A1(_0192_),
    .A2(_0376_),
    .B1(_0378_),
    .Y(_0502_));
 sky130_fd_sc_hd__a221o_1 _1290_ (.A1(_0192_),
    .A2(_0320_),
    .B1(_0374_),
    .B2(_0195_),
    .C1(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__a21oi_1 _1291_ (.A1(_0188_),
    .A2(_0291_),
    .B1(_0289_),
    .Y(_0504_));
 sky130_fd_sc_hd__a221o_1 _1292_ (.A1(_0191_),
    .A2(_0287_),
    .B1(_0278_),
    .B2(_0188_),
    .C1(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__o21ai_1 _1293_ (.A1(_0184_),
    .A2(_0222_),
    .B1(_0224_),
    .Y(_0506_));
 sky130_fd_sc_hd__a221o_1 _1294_ (.A1(_0184_),
    .A2(_0218_),
    .B1(_0220_),
    .B2(_0186_),
    .C1(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__o21ai_1 _1295_ (.A1(_0178_),
    .A2(_0235_),
    .B1(_0237_),
    .Y(_0508_));
 sky130_fd_sc_hd__a221o_1 _1296_ (.A1(_0181_),
    .A2(_0231_),
    .B1(_0232_),
    .B2(_0178_),
    .C1(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__a21oi_1 _1297_ (.A1(\MUL.PS_R1_inst1.LUT_inst14.I1 ),
    .A2(_0240_),
    .B1(_0249_),
    .Y(_0510_));
 sky130_fd_sc_hd__a221oi_4 _1298_ (.A1(\MUL.PS_R1_inst1.LUT_inst13.I1 ),
    .A2(_0242_),
    .B1(_0246_),
    .B2(\MUL.PS_R1_inst1.LUT_inst14.I1 ),
    .C1(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__xnor2_1 _1299_ (.A(_0390_),
    .B(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__xnor2_1 _1300_ (.A(_0509_),
    .B(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__xnor2_1 _1301_ (.A(_0392_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__xnor2_1 _1302_ (.A(_0507_),
    .B(_0514_),
    .Y(_0515_));
 sky130_fd_sc_hd__xnor2_1 _1303_ (.A(_0394_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__xnor2_1 _1304_ (.A(_0505_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__a21oi_1 _1305_ (.A1(_0186_),
    .A2(_0291_),
    .B1(_0289_),
    .Y(_0518_));
 sky130_fd_sc_hd__a221o_1 _1306_ (.A1(_0189_),
    .A2(_0287_),
    .B1(_0278_),
    .B2(_0186_),
    .C1(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__a21oi_1 _1307_ (.A1(\MUL.PS_R1_inst1.LUT_inst15.I1 ),
    .A2(_0248_),
    .B1(_0250_),
    .Y(_0520_));
 sky130_fd_sc_hd__a221o_1 _1308_ (.A1(_0173_),
    .A2(_0243_),
    .B1(_0247_),
    .B2(\MUL.PS_R1_inst1.LUT_inst15.I1 ),
    .C1(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__xor2_2 _1309_ (.A(_0167_),
    .B(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__o21ai_1 _1310_ (.A1(\MUL.PS_R1_inst1.LUT_inst13.I1 ),
    .A2(_0234_),
    .B1(_0236_),
    .Y(_0523_));
 sky130_fd_sc_hd__a221o_1 _1311_ (.A1(_0178_),
    .A2(_0230_),
    .B1(_0232_),
    .B2(_0176_),
    .C1(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__xor2_2 _1312_ (.A(_0511_),
    .B(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__xnor2_1 _1313_ (.A(_0522_),
    .B(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__o21ai_1 _1314_ (.A1(_0181_),
    .A2(_0221_),
    .B1(_0223_),
    .Y(_0527_));
 sky130_fd_sc_hd__a221o_1 _1315_ (.A1(_0181_),
    .A2(_0217_),
    .B1(_0219_),
    .B2(_0184_),
    .C1(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__xnor2_1 _1316_ (.A(_0513_),
    .B(_0528_),
    .Y(_0529_));
 sky130_fd_sc_hd__xnor2_2 _1317_ (.A(_0526_),
    .B(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__xnor2_1 _1318_ (.A(_0515_),
    .B(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__xnor2_2 _1319_ (.A(_0519_),
    .B(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__xor2_1 _1320_ (.A(_0517_),
    .B(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__xnor2_2 _1321_ (.A(_0503_),
    .B(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__o21ai_1 _1322_ (.A1(_0197_),
    .A2(_0402_),
    .B1(_0409_),
    .Y(_0535_));
 sky130_fd_sc_hd__a221o_1 _1323_ (.A1(_0197_),
    .A2(_0423_),
    .B1(_0424_),
    .B2(_0199_),
    .C1(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__a21oi_1 _1324_ (.A1(_0195_),
    .A2(_0376_),
    .B1(_0378_),
    .Y(_0537_));
 sky130_fd_sc_hd__a221o_1 _1325_ (.A1(_0195_),
    .A2(_0319_),
    .B1(_0374_),
    .B2(_0197_),
    .C1(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__xor2_1 _1326_ (.A(_0517_),
    .B(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__xnor2_2 _1327_ (.A(_0398_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__xor2_1 _1328_ (.A(_0536_),
    .B(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__xnor2_2 _1329_ (.A(_0534_),
    .B(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__o21ai_1 _1330_ (.A1(_0199_),
    .A2(_0402_),
    .B1(_0409_),
    .Y(_0543_));
 sky130_fd_sc_hd__a221o_1 _1331_ (.A1(_0199_),
    .A2(_0423_),
    .B1(_0424_),
    .B2(_0201_),
    .C1(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__xnor2_1 _1332_ (.A(_0400_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__xnor2_2 _1333_ (.A(_0540_),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__xor2_1 _1334_ (.A(_0542_),
    .B(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__a21oi_1 _1335_ (.A1(_0501_),
    .A2(_0547_),
    .B1(_0104_),
    .Y(_0548_));
 sky130_fd_sc_hd__o21a_1 _1336_ (.A1(_0501_),
    .A2(_0547_),
    .B1(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__and3_1 _1337_ (.A(\MUL.PS_Rx_inst8.LUT_inst1.i4 ),
    .B(\MUL.PS_Rx_inst8.LUT_inst1.i3 ),
    .C(_0136_),
    .X(_0550_));
 sky130_fd_sc_hd__buf_2 _1338_ (.A(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__a2bb2o_1 _1339_ (.A1_N(_0204_),
    .A2_N(_0498_),
    .B1(_0496_),
    .B2(_0205_),
    .X(_0552_));
 sky130_fd_sc_hd__a211o_1 _1340_ (.A1(_0204_),
    .A2(_0416_),
    .B1(_0551_),
    .C1(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__xnor2_1 _1341_ (.A(_0412_),
    .B(_0546_),
    .Y(_0554_));
 sky130_fd_sc_hd__nand2_1 _1342_ (.A(_0553_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__or2_1 _1343_ (.A(_0553_),
    .B(_0554_),
    .X(_0556_));
 sky130_fd_sc_hd__nand2_2 _1344_ (.A(_0093_),
    .B(_0492_),
    .Y(_0557_));
 sky130_fd_sc_hd__a31o_1 _1345_ (.A1(_0105_),
    .A2(_0555_),
    .A3(_0556_),
    .B1(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__a22oi_1 _1346_ (.A1(_0195_),
    .A2(_0405_),
    .B1(_0424_),
    .B2(_0197_),
    .Y(_0559_));
 sky130_fd_sc_hd__o211a_1 _1347_ (.A1(_0195_),
    .A2(_0402_),
    .B1(_0559_),
    .C1(_0409_),
    .X(_0560_));
 sky130_fd_sc_hd__a21oi_1 _1348_ (.A1(_0188_),
    .A2(_0375_),
    .B1(_0377_),
    .Y(_0561_));
 sky130_fd_sc_hd__a221o_1 _1349_ (.A1(_0189_),
    .A2(_0319_),
    .B1(_0373_),
    .B2(_0192_),
    .C1(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__a21oi_1 _1350_ (.A1(_0184_),
    .A2(_0290_),
    .B1(_0288_),
    .Y(_0563_));
 sky130_fd_sc_hd__a221o_1 _1351_ (.A1(_0186_),
    .A2(_0286_),
    .B1(_0277_),
    .B2(_0184_),
    .C1(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__o21ai_1 _1352_ (.A1(_0178_),
    .A2(_0221_),
    .B1(_0223_),
    .Y(_0565_));
 sky130_fd_sc_hd__a221o_1 _1353_ (.A1(_0178_),
    .A2(_0217_),
    .B1(_0219_),
    .B2(_0181_),
    .C1(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__a21oi_1 _1354_ (.A1(\MUL.PS_R1_inst1.LUT_inst14.I1 ),
    .A2(_0236_),
    .B1(_0234_),
    .Y(_0567_));
 sky130_fd_sc_hd__a221o_1 _1355_ (.A1(_0176_),
    .A2(_0230_),
    .B1(_0232_),
    .B2(\MUL.PS_R1_inst1.LUT_inst14.I1 ),
    .C1(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__inv_2 _1356_ (.A(\MUL.PS_R1_inst1.LUT_inst15.I1 ),
    .Y(_0569_));
 sky130_fd_sc_hd__nand2_1 _1357_ (.A(_0167_),
    .B(\MUL.PS_R1_inst1.LUT_inst14.I1 ),
    .Y(_0570_));
 sky130_fd_sc_hd__o221a_1 _1358_ (.A1(_0167_),
    .A2(_0569_),
    .B1(_0570_),
    .B2(\MUL.PS_Rx_inst2.LUT_inst1.i3 ),
    .C1(_0164_),
    .X(_0571_));
 sky130_fd_sc_hd__a21oi_4 _1359_ (.A1(\MUL.PS_R1_inst1.LUT_inst15.I1 ),
    .A2(_0244_),
    .B1(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__xor2_1 _1360_ (.A(_0568_),
    .B(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__xnor2_1 _1361_ (.A(_0525_),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__xnor2_2 _1362_ (.A(_0566_),
    .B(_0574_),
    .Y(_0575_));
 sky130_fd_sc_hd__xor2_1 _1363_ (.A(_0564_),
    .B(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__xnor2_2 _1364_ (.A(_0530_),
    .B(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__xor2_1 _1365_ (.A(_0562_),
    .B(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__xnor2_1 _1366_ (.A(_0532_),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__xor2_1 _1367_ (.A(_0560_),
    .B(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__xnor2_2 _1368_ (.A(_0534_),
    .B(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__a2bb2o_1 _1369_ (.A1_N(_0199_),
    .A2_N(_0498_),
    .B1(_0496_),
    .B2(_0202_),
    .X(_0582_));
 sky130_fd_sc_hd__a211o_1 _1370_ (.A1(_0199_),
    .A2(_0416_),
    .B1(_0551_),
    .C1(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__xor2_1 _1371_ (.A(_0581_),
    .B(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__nand2_1 _1372_ (.A(_0542_),
    .B(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__o21a_1 _1373_ (.A1(_0542_),
    .A2(_0584_),
    .B1(_0104_),
    .X(_0586_));
 sky130_fd_sc_hd__a2bb2o_1 _1374_ (.A1_N(_0197_),
    .A2_N(_0497_),
    .B1(_0495_),
    .B2(_0199_),
    .X(_0587_));
 sky130_fd_sc_hd__a211o_1 _1375_ (.A1(_0197_),
    .A2(_0415_),
    .B1(_0551_),
    .C1(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__o21ai_1 _1376_ (.A1(_0169_),
    .A2(_0235_),
    .B1(_0237_),
    .Y(_0589_));
 sky130_fd_sc_hd__a221o_1 _1377_ (.A1(_0173_),
    .A2(_0231_),
    .B1(_0233_),
    .B2(_0169_),
    .C1(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__xnor2_2 _1378_ (.A(_0479_),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__xnor2_4 _1379_ (.A(_0572_),
    .B(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__xnor2_1 _1380_ (.A(_0522_),
    .B(_0573_),
    .Y(_0593_));
 sky130_fd_sc_hd__o21ai_1 _1381_ (.A1(_0176_),
    .A2(_0222_),
    .B1(_0224_),
    .Y(_0594_));
 sky130_fd_sc_hd__a221o_1 _1382_ (.A1(_0176_),
    .A2(_0218_),
    .B1(_0220_),
    .B2(_0178_),
    .C1(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__xnor2_2 _1383_ (.A(_0593_),
    .B(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__xnor2_4 _1384_ (.A(_0592_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__a21oi_1 _1385_ (.A1(_0181_),
    .A2(_0291_),
    .B1(_0289_),
    .Y(_0598_));
 sky130_fd_sc_hd__a221o_1 _1386_ (.A1(_0184_),
    .A2(_0287_),
    .B1(_0278_),
    .B2(_0181_),
    .C1(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__xor2_1 _1387_ (.A(_0575_),
    .B(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__xnor2_2 _1388_ (.A(_0597_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__xnor2_1 _1389_ (.A(_0577_),
    .B(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__a21oi_1 _1390_ (.A1(_0187_),
    .A2(_0376_),
    .B1(_0378_),
    .Y(_0603_));
 sky130_fd_sc_hd__a221o_1 _1391_ (.A1(_0187_),
    .A2(_0320_),
    .B1(_0374_),
    .B2(_0189_),
    .C1(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__xnor2_2 _1392_ (.A(_0602_),
    .B(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__o21ai_1 _1393_ (.A1(_0192_),
    .A2(_0401_),
    .B1(_0408_),
    .Y(_0606_));
 sky130_fd_sc_hd__a221o_1 _1394_ (.A1(_0192_),
    .A2(_0423_),
    .B1(_0424_),
    .B2(_0195_),
    .C1(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__xnor2_1 _1395_ (.A(_0579_),
    .B(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__xnor2_2 _1396_ (.A(_0605_),
    .B(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__xnor2_1 _1397_ (.A(_0588_),
    .B(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__a21oi_1 _1398_ (.A1(_0581_),
    .A2(_0610_),
    .B1(_0104_),
    .Y(_0611_));
 sky130_fd_sc_hd__o21a_1 _1399_ (.A1(_0581_),
    .A2(_0610_),
    .B1(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__a211o_1 _1400_ (.A1(_0585_),
    .A2(_0586_),
    .B1(_0102_),
    .C1(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__o21a_1 _1401_ (.A1(_0549_),
    .A2(_0558_),
    .B1(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__a21oi_1 _1402_ (.A1(_0185_),
    .A2(_0376_),
    .B1(_0378_),
    .Y(_0615_));
 sky130_fd_sc_hd__a221o_1 _1403_ (.A1(_0185_),
    .A2(_0320_),
    .B1(_0374_),
    .B2(_0187_),
    .C1(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__xor2_2 _1404_ (.A(_0601_),
    .B(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__and2_1 _1405_ (.A(_0173_),
    .B(_0224_),
    .X(_0618_));
 sky130_fd_sc_hd__nor2_1 _1406_ (.A(_0222_),
    .B(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__a221o_1 _1407_ (.A1(_0173_),
    .A2(_0218_),
    .B1(_0220_),
    .B2(_0176_),
    .C1(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__xor2_2 _1408_ (.A(_0592_),
    .B(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__a21oi_1 _1409_ (.A1(_0178_),
    .A2(_0291_),
    .B1(_0289_),
    .Y(_0622_));
 sky130_fd_sc_hd__a221o_1 _1410_ (.A1(_0181_),
    .A2(_0287_),
    .B1(_0278_),
    .B2(_0178_),
    .C1(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__nor2_1 _1411_ (.A(_0160_),
    .B(_0169_),
    .Y(_0624_));
 sky130_fd_sc_hd__a2bb2oi_1 _1412_ (.A1_N(_0164_),
    .A2_N(_0169_),
    .B1(_0228_),
    .B2(_0227_),
    .Y(_0625_));
 sky130_fd_sc_hd__inv_2 _1413_ (.A(_0173_),
    .Y(_0626_));
 sky130_fd_sc_hd__o211a_1 _1414_ (.A1(\MUL.PS_Rx_inst3.LUT_inst1.i3 ),
    .A2(_0626_),
    .B1(_0164_),
    .C1(_0160_),
    .X(_0627_));
 sky130_fd_sc_hd__o21ba_1 _1415_ (.A1(_0624_),
    .A2(_0625_),
    .B1_N(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__xnor2_1 _1416_ (.A(_0623_),
    .B(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__xnor2_1 _1417_ (.A(_0621_),
    .B(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__xnor2_2 _1418_ (.A(_0597_),
    .B(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__o21ai_1 _1419_ (.A1(_0189_),
    .A2(_0401_),
    .B1(_0409_),
    .Y(_0632_));
 sky130_fd_sc_hd__a221o_1 _1420_ (.A1(_0189_),
    .A2(_0423_),
    .B1(_0424_),
    .B2(_0192_),
    .C1(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__xnor2_1 _1421_ (.A(_0631_),
    .B(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__xnor2_1 _1422_ (.A(_0617_),
    .B(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__xnor2_2 _1423_ (.A(_0605_),
    .B(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__a2bb2o_1 _1424_ (.A1_N(_0195_),
    .A2_N(_0498_),
    .B1(_0496_),
    .B2(_0197_),
    .X(_0637_));
 sky130_fd_sc_hd__a211o_1 _1425_ (.A1(_0195_),
    .A2(_0416_),
    .B1(_0551_),
    .C1(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__xnor2_1 _1426_ (.A(_0636_),
    .B(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__a21boi_1 _1427_ (.A1(_0609_),
    .A2(_0639_),
    .B1_N(_0104_),
    .Y(_0640_));
 sky130_fd_sc_hd__o21ai_1 _1428_ (.A1(_0609_),
    .A2(_0639_),
    .B1(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__a2bb2o_1 _1429_ (.A1_N(_0192_),
    .A2_N(_0498_),
    .B1(_0496_),
    .B2(_0195_),
    .X(_0642_));
 sky130_fd_sc_hd__a211o_1 _1430_ (.A1(_0192_),
    .A2(_0416_),
    .B1(_0551_),
    .C1(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__a21oi_1 _1431_ (.A1(_0182_),
    .A2(_0375_),
    .B1(_0377_),
    .Y(_0644_));
 sky130_fd_sc_hd__a221o_1 _1432_ (.A1(_0182_),
    .A2(_0319_),
    .B1(_0373_),
    .B2(_0185_),
    .C1(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__o21ai_1 _1433_ (.A1(_0169_),
    .A2(_0222_),
    .B1(_0224_),
    .Y(_0646_));
 sky130_fd_sc_hd__a221o_1 _1434_ (.A1(_0169_),
    .A2(_0218_),
    .B1(_0220_),
    .B2(_0173_),
    .C1(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__xnor2_2 _1435_ (.A(_0479_),
    .B(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__a21oi_1 _1436_ (.A1(_0176_),
    .A2(_0291_),
    .B1(_0289_),
    .Y(_0649_));
 sky130_fd_sc_hd__a221o_1 _1437_ (.A1(_0178_),
    .A2(_0287_),
    .B1(_0278_),
    .B2(_0176_),
    .C1(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__xnor2_1 _1438_ (.A(_0648_),
    .B(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__xnor2_2 _1439_ (.A(_0621_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__xnor2_1 _1440_ (.A(_0645_),
    .B(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__o21ai_1 _1441_ (.A1(_0187_),
    .A2(_0401_),
    .B1(_0408_),
    .Y(_0654_));
 sky130_fd_sc_hd__a221o_1 _1442_ (.A1(_0187_),
    .A2(_0405_),
    .B1(_0406_),
    .B2(_0189_),
    .C1(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__xnor2_1 _1443_ (.A(_0653_),
    .B(_0655_),
    .Y(_0656_));
 sky130_fd_sc_hd__xnor2_2 _1444_ (.A(_0617_),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__xor2_1 _1445_ (.A(_0643_),
    .B(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__a21oi_1 _1446_ (.A1(_0636_),
    .A2(_0658_),
    .B1(_0105_),
    .Y(_0659_));
 sky130_fd_sc_hd__o21ai_1 _1447_ (.A1(_0636_),
    .A2(_0658_),
    .B1(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__nor2_1 _1448_ (.A(_0153_),
    .B(_0169_),
    .Y(_0661_));
 sky130_fd_sc_hd__o21ba_1 _1449_ (.A1(_0153_),
    .A2(_0216_),
    .B1_N(_0624_),
    .X(_0662_));
 sky130_fd_sc_hd__o32a_1 _1450_ (.A1(_0279_),
    .A2(_0227_),
    .A3(_0618_),
    .B1(_0661_),
    .B2(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__xnor2_1 _1451_ (.A(_0628_),
    .B(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__and2_1 _1452_ (.A(_0173_),
    .B(_0290_),
    .X(_0665_));
 sky130_fd_sc_hd__nor2_1 _1453_ (.A(_0289_),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__a221o_1 _1454_ (.A1(_0176_),
    .A2(_0287_),
    .B1(_0277_),
    .B2(_0173_),
    .C1(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__xnor2_1 _1455_ (.A(_0664_),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__xnor2_2 _1456_ (.A(_0648_),
    .B(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__a21oi_1 _1457_ (.A1(_0179_),
    .A2(_0376_),
    .B1(_0378_),
    .Y(_0670_));
 sky130_fd_sc_hd__a221o_1 _1458_ (.A1(_0179_),
    .A2(_0320_),
    .B1(_0374_),
    .B2(_0182_),
    .C1(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__xnor2_1 _1459_ (.A(_0669_),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__xnor2_1 _1460_ (.A(_0645_),
    .B(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__o21ai_1 _1461_ (.A1(_0185_),
    .A2(_0402_),
    .B1(_0409_),
    .Y(_0674_));
 sky130_fd_sc_hd__a221o_1 _1462_ (.A1(_0185_),
    .A2(_0423_),
    .B1(_0424_),
    .B2(_0187_),
    .C1(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__xnor2_1 _1463_ (.A(_0631_),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__xnor2_1 _1464_ (.A(_0673_),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__a2bb2o_1 _1465_ (.A1_N(_0187_),
    .A2_N(_0497_),
    .B1(_0495_),
    .B2(_0189_),
    .X(_0678_));
 sky130_fd_sc_hd__a211o_1 _1466_ (.A1(_0187_),
    .A2(_0415_),
    .B1(_0550_),
    .C1(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__xnor2_1 _1467_ (.A(_0652_),
    .B(_0672_),
    .Y(_0680_));
 sky130_fd_sc_hd__a21oi_1 _1468_ (.A1(_0177_),
    .A2(_0375_),
    .B1(_0377_),
    .Y(_0681_));
 sky130_fd_sc_hd__a221o_1 _1469_ (.A1(_0177_),
    .A2(_0319_),
    .B1(_0373_),
    .B2(_0179_),
    .C1(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__a21oi_1 _1470_ (.A1(_0169_),
    .A2(_0290_),
    .B1(_0288_),
    .Y(_0683_));
 sky130_fd_sc_hd__a221o_1 _1471_ (.A1(_0173_),
    .A2(_0286_),
    .B1(_0277_),
    .B2(_0169_),
    .C1(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__xnor2_1 _1472_ (.A(_0478_),
    .B(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__xnor2_2 _1473_ (.A(_0663_),
    .B(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__xor2_1 _1474_ (.A(_0682_),
    .B(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__xnor2_2 _1475_ (.A(_0669_),
    .B(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__o21ai_1 _1476_ (.A1(_0182_),
    .A2(_0401_),
    .B1(_0408_),
    .Y(_0689_));
 sky130_fd_sc_hd__a221o_1 _1477_ (.A1(_0182_),
    .A2(_0405_),
    .B1(_0406_),
    .B2(_0185_),
    .C1(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__xnor2_1 _1478_ (.A(_0688_),
    .B(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__xnor2_2 _1479_ (.A(_0680_),
    .B(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__xor2_1 _1480_ (.A(_0679_),
    .B(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__a2bb2o_1 _1481_ (.A1_N(_0189_),
    .A2_N(_0497_),
    .B1(_0495_),
    .B2(_0192_),
    .X(_0694_));
 sky130_fd_sc_hd__a211o_1 _1482_ (.A1(_0189_),
    .A2(_0415_),
    .B1(_0550_),
    .C1(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__xnor2_1 _1483_ (.A(_0657_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__mux2_1 _1484_ (.A0(_0693_),
    .A1(_0696_),
    .S(\count2[0] ),
    .X(_0697_));
 sky130_fd_sc_hd__xnor2_1 _1485_ (.A(_0677_),
    .B(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__o21ai_1 _1486_ (.A1(_0102_),
    .A2(_0698_),
    .B1(_0494_),
    .Y(_0699_));
 sky130_fd_sc_hd__a31o_1 _1487_ (.A1(_0102_),
    .A2(_0641_),
    .A3(_0660_),
    .B1(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__or2_1 _1488_ (.A(\count2[3] ),
    .B(_0491_),
    .X(_0701_));
 sky130_fd_sc_hd__nand3_1 _1489_ (.A(\count2[5] ),
    .B(\count2[4] ),
    .C(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__nand2_1 _1490_ (.A(\count2[3] ),
    .B(_0491_),
    .Y(_0703_));
 sky130_fd_sc_hd__and2_1 _1491_ (.A(_0701_),
    .B(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__o2111a_1 _1492_ (.A1(_0494_),
    .A2(_0614_),
    .B1(_0700_),
    .C1(_0702_),
    .D1(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__a21oi_1 _1493_ (.A1(_0170_),
    .A2(_0376_),
    .B1(_0378_),
    .Y(_0706_));
 sky130_fd_sc_hd__a221o_1 _1494_ (.A1(_0170_),
    .A2(_0320_),
    .B1(_0374_),
    .B2(_0174_),
    .C1(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__nor2_1 _1495_ (.A(_0150_),
    .B(_0170_),
    .Y(_0708_));
 sky130_fd_sc_hd__o21ba_1 _1496_ (.A1(_0150_),
    .A2(_0276_),
    .B1_N(_0661_),
    .X(_0709_));
 sky130_fd_sc_hd__o32a_1 _1497_ (.A1(_0321_),
    .A2(_0279_),
    .A3(_0665_),
    .B1(_0708_),
    .B2(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__xnor2_1 _1498_ (.A(_0478_),
    .B(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__xnor2_2 _1499_ (.A(_0707_),
    .B(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__o211a_1 _1500_ (.A1(\MUL.PS_Rx_inst6.LUT_inst1.i3 ),
    .A2(_0626_),
    .B1(_0150_),
    .C1(_0141_),
    .X(_0713_));
 sky130_fd_sc_hd__a221o_1 _1501_ (.A1(_0170_),
    .A2(_0318_),
    .B1(_0708_),
    .B2(_0141_),
    .C1(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__and2_1 _1502_ (.A(_0174_),
    .B(_0408_),
    .X(_0715_));
 sky130_fd_sc_hd__nor2_1 _1503_ (.A(_0402_),
    .B(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__a221o_1 _1504_ (.A1(_0174_),
    .A2(_0423_),
    .B1(_0424_),
    .B2(_0177_),
    .C1(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__xnor2_1 _1505_ (.A(_0714_),
    .B(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__xnor2_2 _1506_ (.A(_0712_),
    .B(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__a21oi_1 _1507_ (.A1(_0170_),
    .A2(_0409_),
    .B1(_0402_),
    .Y(_0720_));
 sky130_fd_sc_hd__a221o_1 _1508_ (.A1(_0170_),
    .A2(_0423_),
    .B1(_0424_),
    .B2(_0174_),
    .C1(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__xnor2_1 _1509_ (.A(_0479_),
    .B(_0714_),
    .Y(_0722_));
 sky130_fd_sc_hd__xnor2_2 _1510_ (.A(_0721_),
    .B(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__a2bb2o_1 _1511_ (.A1_N(_0177_),
    .A2_N(_0497_),
    .B1(_0495_),
    .B2(_0179_),
    .X(_0724_));
 sky130_fd_sc_hd__a211o_1 _1512_ (.A1(_0177_),
    .A2(_0415_),
    .B1(_0551_),
    .C1(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__xnor2_1 _1513_ (.A(_0723_),
    .B(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__nand2_1 _1514_ (.A(_0719_),
    .B(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__or2_1 _1515_ (.A(_0719_),
    .B(_0726_),
    .X(_0728_));
 sky130_fd_sc_hd__a21oi_1 _1516_ (.A1(_0174_),
    .A2(_0375_),
    .B1(_0377_),
    .Y(_0729_));
 sky130_fd_sc_hd__a221o_1 _1517_ (.A1(_0174_),
    .A2(_0319_),
    .B1(_0373_),
    .B2(_0177_),
    .C1(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__xor2_1 _1518_ (.A(_0710_),
    .B(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__xnor2_2 _1519_ (.A(_0686_),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__o21ai_1 _1520_ (.A1(_0179_),
    .A2(_0402_),
    .B1(_0409_),
    .Y(_0733_));
 sky130_fd_sc_hd__a221o_1 _1521_ (.A1(_0179_),
    .A2(_0423_),
    .B1(_0424_),
    .B2(_0182_),
    .C1(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__xor2_1 _1522_ (.A(_0732_),
    .B(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__xnor2_2 _1523_ (.A(_0688_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__a22oi_1 _1524_ (.A1(_0177_),
    .A2(_0405_),
    .B1(_0406_),
    .B2(_0179_),
    .Y(_0737_));
 sky130_fd_sc_hd__o211a_1 _1525_ (.A1(_0177_),
    .A2(_0402_),
    .B1(_0737_),
    .C1(_0409_),
    .X(_0738_));
 sky130_fd_sc_hd__xnor2_1 _1526_ (.A(_0712_),
    .B(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__xnor2_2 _1527_ (.A(_0732_),
    .B(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__a2bb2o_1 _1528_ (.A1_N(_0182_),
    .A2_N(_0498_),
    .B1(_0496_),
    .B2(_0185_),
    .X(_0741_));
 sky130_fd_sc_hd__a211o_1 _1529_ (.A1(_0182_),
    .A2(_0416_),
    .B1(_0551_),
    .C1(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__xnor2_1 _1530_ (.A(_0740_),
    .B(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__or2_1 _1531_ (.A(_0736_),
    .B(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__a21oi_1 _1532_ (.A1(_0736_),
    .A2(_0743_),
    .B1(_0332_),
    .Y(_0745_));
 sky130_fd_sc_hd__a32o_1 _1533_ (.A1(_0332_),
    .A2(_0727_),
    .A3(_0728_),
    .B1(_0744_),
    .B2(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__a2bb2o_1 _1534_ (.A1_N(_0179_),
    .A2_N(_0498_),
    .B1(_0496_),
    .B2(_0182_),
    .X(_0747_));
 sky130_fd_sc_hd__a211o_1 _1535_ (.A1(_0179_),
    .A2(_0416_),
    .B1(_0551_),
    .C1(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__xor2_1 _1536_ (.A(_0719_),
    .B(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__nand2_1 _1537_ (.A(_0740_),
    .B(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__o21a_1 _1538_ (.A1(_0740_),
    .A2(_0749_),
    .B1(\count2[1] ),
    .X(_0751_));
 sky130_fd_sc_hd__a2bb2o_1 _1539_ (.A1_N(_0185_),
    .A2_N(_0498_),
    .B1(_0496_),
    .B2(_0187_),
    .X(_0752_));
 sky130_fd_sc_hd__a211o_1 _1540_ (.A1(_0185_),
    .A2(_0416_),
    .B1(_0551_),
    .C1(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__xor2_1 _1541_ (.A(_0736_),
    .B(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__or2_1 _1542_ (.A(_0692_),
    .B(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__a21oi_1 _1543_ (.A1(_0692_),
    .A2(_0754_),
    .B1(_0557_),
    .Y(_0756_));
 sky130_fd_sc_hd__a22o_1 _1544_ (.A1(_0750_),
    .A2(_0751_),
    .B1(_0755_),
    .B2(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_1 _1545_ (.A0(_0746_),
    .A1(_0757_),
    .S(_0105_),
    .X(_0758_));
 sky130_fd_sc_hd__nor2_1 _1546_ (.A(_0136_),
    .B(_0170_),
    .Y(_0759_));
 sky130_fd_sc_hd__o22a_1 _1547_ (.A1(_0141_),
    .A2(_0170_),
    .B1(_0404_),
    .B2(_0136_),
    .X(_0760_));
 sky130_fd_sc_hd__o32a_1 _1548_ (.A1(_0417_),
    .A2(_0443_),
    .A3(_0715_),
    .B1(_0759_),
    .B2(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__or3_1 _1549_ (.A(\MUL.PS_Rx_inst8.LUT_inst1.i4 ),
    .B(_0569_),
    .C(_0414_),
    .X(_0762_));
 sky130_fd_sc_hd__o2bb2a_1 _1550_ (.A1_N(_0174_),
    .A2_N(_0496_),
    .B1(_0762_),
    .B2(_0413_),
    .X(_0763_));
 sky130_fd_sc_hd__o211a_1 _1551_ (.A1(_0170_),
    .A2(_0498_),
    .B1(_0499_),
    .C1(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__xnor2_1 _1552_ (.A(_0478_),
    .B(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__and2_1 _1553_ (.A(_0761_),
    .B(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__nor2_1 _1554_ (.A(_0761_),
    .B(_0765_),
    .Y(_0767_));
 sky130_fd_sc_hd__a21oi_1 _1555_ (.A1(_0174_),
    .A2(_0499_),
    .B1(_0498_),
    .Y(_0768_));
 sky130_fd_sc_hd__a221o_1 _1556_ (.A1(_0174_),
    .A2(_0416_),
    .B1(_0496_),
    .B2(_0177_),
    .C1(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__xor2_1 _1557_ (.A(_0769_),
    .B(_0761_),
    .X(_0770_));
 sky130_fd_sc_hd__nor2_1 _1558_ (.A(_0723_),
    .B(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__a21bo_1 _1559_ (.A1(_0723_),
    .A2(_0770_),
    .B1_N(_0104_),
    .X(_0772_));
 sky130_fd_sc_hd__o32a_1 _1560_ (.A1(_0105_),
    .A2(_0766_),
    .A3(_0767_),
    .B1(_0771_),
    .B2(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__o21a_1 _1561_ (.A1(_0626_),
    .A2(_0551_),
    .B1(_0136_),
    .X(_0774_));
 sky130_fd_sc_hd__o21ai_1 _1562_ (.A1(_0759_),
    .A2(_0774_),
    .B1(\MUL.PS_Rx_inst8.LUT_inst1.i4 ),
    .Y(_0775_));
 sky130_fd_sc_hd__a32o_1 _1563_ (.A1(_0094_),
    .A2(_0762_),
    .A3(_0775_),
    .B1(_0479_),
    .B2(_0493_),
    .X(_0776_));
 sky130_fd_sc_hd__and2_1 _1564_ (.A(_0491_),
    .B(_0493_),
    .X(_0777_));
 sky130_fd_sc_hd__a211o_1 _1565_ (.A1(_0102_),
    .A2(_0773_),
    .B1(_0776_),
    .C1(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__nand2_1 _1566_ (.A(_0701_),
    .B(_0703_),
    .Y(_0779_));
 sky130_fd_sc_hd__o2111a_1 _1567_ (.A1(_0494_),
    .A2(_0758_),
    .B1(_0778_),
    .C1(_0702_),
    .D1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__xnor2_1 _1568_ (.A(\count2[4] ),
    .B(_0701_),
    .Y(_0781_));
 sky130_fd_sc_hd__o21ba_1 _1569_ (.A1(_0705_),
    .A2(_0780_),
    .B1_N(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__nor2_1 _1570_ (.A(_0492_),
    .B(_0422_),
    .Y(_0783_));
 sky130_fd_sc_hd__nor2_1 _1571_ (.A(_0093_),
    .B(_0436_),
    .Y(_0784_));
 sky130_fd_sc_hd__a221o_1 _1572_ (.A1(_0464_),
    .A2(_0448_),
    .B1(_0449_),
    .B2(_0440_),
    .C1(_0777_),
    .X(_0785_));
 sky130_fd_sc_hd__or3_1 _1573_ (.A(_0783_),
    .B(_0784_),
    .C(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__nor2_1 _1574_ (.A(_0492_),
    .B(_0326_),
    .Y(_0787_));
 sky130_fd_sc_hd__mux2_1 _1575_ (.A0(_0284_),
    .A1(_0264_),
    .S(_0104_),
    .X(_0788_));
 sky130_fd_sc_hd__o21ai_1 _1576_ (.A1(_0557_),
    .A2(_0788_),
    .B1(_0777_),
    .Y(_0789_));
 sky130_fd_sc_hd__a211o_1 _1577_ (.A1(_0094_),
    .A2(_0330_),
    .B1(_0787_),
    .C1(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__mux4_1 _1578_ (.A0(_0457_),
    .A1(_0463_),
    .A2(_0484_),
    .A3(_0476_),
    .S0(_0104_),
    .S1(_0777_),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _1579_ (.A0(_0469_),
    .A1(_0471_),
    .S(_0104_),
    .X(_0792_));
 sky130_fd_sc_hd__mux2_1 _1580_ (.A0(_0486_),
    .A1(_0206_),
    .S(\count2[0] ),
    .X(_0793_));
 sky130_fd_sc_hd__a21o_1 _1581_ (.A1(_0777_),
    .A2(_0793_),
    .B1(_0557_),
    .X(_0794_));
 sky130_fd_sc_hd__a21o_1 _1582_ (.A1(_0494_),
    .A2(_0792_),
    .B1(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__o211a_1 _1583_ (.A1(_0102_),
    .A2(_0791_),
    .B1(_0795_),
    .C1(_0704_),
    .X(_0796_));
 sky130_fd_sc_hd__a31o_1 _1584_ (.A1(_0779_),
    .A2(_0786_),
    .A3(_0790_),
    .B1(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__a311o_1 _1585_ (.A1(_0781_),
    .A2(_0702_),
    .A3(_0797_),
    .B1(_0098_),
    .C1(_0209_),
    .X(_0798_));
 sky130_fd_sc_hd__o22a_1 _1586_ (.A1(net7),
    .A2(_0214_),
    .B1(_0782_),
    .B2(_0798_),
    .X(_0077_));
 sky130_fd_sc_hd__inv_2 _1587_ (.A(_0213_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _1588_ (.A(_0213_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1589_ (.A(_0213_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _1590_ (.A(_0213_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1591_ (.A(_0213_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _1592_ (.A(_0213_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _1593_ (.A(_0213_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _1594_ (.A(_0213_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1595_ (.A(_0209_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _1596_ (.A(_0209_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _1597_ (.A(_0209_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _1598_ (.A(_0209_),
    .Y(_0043_));
 sky130_fd_sc_hd__dfrtp_1 _1599_ (.CLK(net11),
    .D(_0044_),
    .RESET_B(_0000_),
    .Q(\MUL.PS_R1_inst1.LUT_inst1.i0 ));
 sky130_fd_sc_hd__dfrtp_4 _1600_ (.CLK(net10),
    .D(_0045_),
    .RESET_B(_0001_),
    .Q(\MUL.PS_R1_inst1.LUT_inst1.i1 ));
 sky130_fd_sc_hd__dfrtp_2 _1601_ (.CLK(clknet_1_1__leaf_net8),
    .D(_0046_),
    .RESET_B(_0002_),
    .Q(\MUL.PS_R1_inst1.LUT_inst2.I1 ));
 sky130_fd_sc_hd__dfrtp_2 _1602_ (.CLK(net13),
    .D(_0047_),
    .RESET_B(_0003_),
    .Q(\MUL.PS_R1_inst1.LUT_inst3.I1 ));
 sky130_fd_sc_hd__dfrtp_1 _1603_ (.CLK(net9),
    .D(_0048_),
    .RESET_B(_0004_),
    .Q(\MUL.PS_R1_inst1.LUT_inst4.I1 ));
 sky130_fd_sc_hd__dfrtp_4 _1604_ (.CLK(net10),
    .D(_0049_),
    .RESET_B(_0005_),
    .Q(\MUL.PS_R1_inst1.LUT_inst5.I1 ));
 sky130_fd_sc_hd__dfrtp_2 _1605_ (.CLK(clknet_1_1__leaf_net8),
    .D(_0050_),
    .RESET_B(_0006_),
    .Q(\MUL.PS_R1_inst1.LUT_inst6.I1 ));
 sky130_fd_sc_hd__dfrtp_2 _1606_ (.CLK(net9),
    .D(_0051_),
    .RESET_B(_0007_),
    .Q(\MUL.PS_R1_inst1.LUT_inst7.I1 ));
 sky130_fd_sc_hd__dfrtp_4 _1607_ (.CLK(clknet_1_0__leaf_net8),
    .D(_0052_),
    .RESET_B(_0008_),
    .Q(\MUL.PS_R1_inst1.LUT_inst8.I1 ));
 sky130_fd_sc_hd__dfrtp_2 _1608_ (.CLK(net9),
    .D(_0053_),
    .RESET_B(_0009_),
    .Q(\MUL.PS_R1_inst1.LUT_inst10.I0 ));
 sky130_fd_sc_hd__dfrtp_2 _1609_ (.CLK(clknet_1_1__leaf_net8),
    .D(_0054_),
    .RESET_B(_0010_),
    .Q(\MUL.PS_R1_inst1.LUT_inst10.I1 ));
 sky130_fd_sc_hd__dfrtp_4 _1610_ (.CLK(net9),
    .D(_0055_),
    .RESET_B(_0011_),
    .Q(\MUL.PS_R1_inst1.LUT_inst11.I1 ));
 sky130_fd_sc_hd__dfrtp_4 _1611_ (.CLK(net9),
    .D(_0056_),
    .RESET_B(_0012_),
    .Q(\MUL.PS_R1_inst1.LUT_inst12.I1 ));
 sky130_fd_sc_hd__dfrtp_2 _1612_ (.CLK(net9),
    .D(_0057_),
    .RESET_B(_0013_),
    .Q(\MUL.PS_R1_inst1.LUT_inst13.I1 ));
 sky130_fd_sc_hd__dfrtp_4 _1613_ (.CLK(clknet_1_1__leaf_net8),
    .D(_0058_),
    .RESET_B(_0014_),
    .Q(\MUL.PS_R1_inst1.LUT_inst14.I1 ));
 sky130_fd_sc_hd__dfrtp_4 _1614_ (.CLK(net13),
    .D(_0059_),
    .RESET_B(_0015_),
    .Q(\MUL.PS_R1_inst1.LUT_inst15.I1 ));
 sky130_fd_sc_hd__dfrtp_1 _1615_ (.CLK(net10),
    .D(_0060_),
    .RESET_B(_0016_),
    .Q(\MUL.PS_R1_inst1.LUT_inst1.i3 ));
 sky130_fd_sc_hd__dfrtp_1 _1616_ (.CLK(net9),
    .D(_0061_),
    .RESET_B(_0017_),
    .Q(\MUL.PS_R1_inst1.LUT_inst1.i4 ));
 sky130_fd_sc_hd__dfrtp_2 _1617_ (.CLK(clknet_1_0__leaf_net8),
    .D(_0062_),
    .RESET_B(_0018_),
    .Q(\MUL.PS_Rx_inst2.LUT_inst1.i3 ));
 sky130_fd_sc_hd__dfrtp_1 _1618_ (.CLK(net9),
    .D(_0063_),
    .RESET_B(_0019_),
    .Q(\MUL.PS_Rx_inst2.LUT_inst1.i4 ));
 sky130_fd_sc_hd__dfrtp_2 _1619_ (.CLK(clknet_1_1__leaf_net8),
    .D(_0064_),
    .RESET_B(_0020_),
    .Q(\MUL.PS_Rx_inst3.LUT_inst1.i3 ));
 sky130_fd_sc_hd__dfrtp_1 _1620_ (.CLK(net9),
    .D(_0065_),
    .RESET_B(_0021_),
    .Q(\MUL.PS_Rx_inst3.LUT_inst1.i4 ));
 sky130_fd_sc_hd__dfrtp_2 _1621_ (.CLK(clknet_1_1__leaf_net8),
    .D(_0066_),
    .RESET_B(_0022_),
    .Q(\MUL.PS_Rx_inst4.LUT_inst1.i3 ));
 sky130_fd_sc_hd__dfrtp_1 _1622_ (.CLK(net9),
    .D(_0067_),
    .RESET_B(_0023_),
    .Q(\MUL.PS_Rx_inst4.LUT_inst1.i4 ));
 sky130_fd_sc_hd__dfrtp_4 _1623_ (.CLK(clknet_1_0__leaf_net8),
    .D(_0068_),
    .RESET_B(_0024_),
    .Q(\MUL.PS_Rx_inst5.LUT_inst1.i3 ));
 sky130_fd_sc_hd__dfrtp_2 _1624_ (.CLK(net13),
    .D(_0069_),
    .RESET_B(_0025_),
    .Q(\MUL.PS_Rx_inst5.LUT_inst1.i4 ));
 sky130_fd_sc_hd__dfrtp_4 _1625_ (.CLK(net11),
    .D(_0070_),
    .RESET_B(_0026_),
    .Q(\MUL.PS_Rx_inst6.LUT_inst1.i3 ));
 sky130_fd_sc_hd__dfrtp_2 _1626_ (.CLK(net13),
    .D(_0071_),
    .RESET_B(_0027_),
    .Q(\MUL.PS_Rx_inst6.LUT_inst1.i4 ));
 sky130_fd_sc_hd__dfrtp_2 _1627_ (.CLK(net11),
    .D(_0072_),
    .RESET_B(_0028_),
    .Q(\MUL.PS_Rx_inst7.LUT_inst1.i3 ));
 sky130_fd_sc_hd__dfrtp_4 _1628_ (.CLK(net11),
    .D(_0073_),
    .RESET_B(_0029_),
    .Q(\MUL.PS_Rx_inst7.LUT_inst1.i4 ));
 sky130_fd_sc_hd__dfrtp_2 _1629_ (.CLK(net11),
    .D(_0074_),
    .RESET_B(_0030_),
    .Q(\MUL.PS_Rx_inst8.LUT_inst1.i3 ));
 sky130_fd_sc_hd__dfrtp_4 _1630_ (.CLK(net11),
    .D(_0075_),
    .RESET_B(_0031_),
    .Q(\MUL.PS_Rx_inst8.LUT_inst1.i4 ));
 sky130_fd_sc_hd__dfxtp_1 _1631_ (.CLK(clknet_1_1__leaf_net12),
    .D(_0076_),
    .Q(net6));
 sky130_fd_sc_hd__dfxtp_2 _1632_ (.CLK(clknet_1_1__leaf_net12),
    .D(_0077_),
    .Q(net7));
 sky130_fd_sc_hd__dfrtp_2 _1633_ (.CLK(net10),
    .D(_0078_),
    .RESET_B(_0032_),
    .Q(\count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1634_ (.CLK(clknet_1_0__leaf_net8),
    .D(_0079_),
    .RESET_B(_0033_),
    .Q(\count[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1635_ (.CLK(net11),
    .D(_0080_),
    .RESET_B(_0034_),
    .Q(\count[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1636_ (.CLK(net11),
    .D(_0081_),
    .RESET_B(_0035_),
    .Q(\count[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1637_ (.CLK(net10),
    .D(_0082_),
    .RESET_B(_0036_),
    .Q(\count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1638_ (.CLK(net10),
    .D(_0083_),
    .RESET_B(_0037_),
    .Q(\count[5] ));
 sky130_fd_sc_hd__dfrtp_4 _1639_ (.CLK(net11),
    .D(_0084_),
    .RESET_B(_0038_),
    .Q(\count2[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1640_ (.CLK(net11),
    .D(_0085_),
    .RESET_B(_0039_),
    .Q(\count2[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1641_ (.CLK(clknet_1_1__leaf_net12),
    .D(_0086_),
    .RESET_B(_0040_),
    .Q(\count2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1642_ (.CLK(clknet_1_0__leaf_net12),
    .D(_0087_),
    .RESET_B(_0041_),
    .Q(\count2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1643_ (.CLK(clknet_1_0__leaf_net12),
    .D(_0088_),
    .RESET_B(_0042_),
    .Q(\count2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1644_ (.CLK(clknet_1_0__leaf_net12),
    .D(_0089_),
    .RESET_B(_0043_),
    .Q(\count2[5] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(A_PAD),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(B_PAD),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(sel),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(user_clock2),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(wb_rst_i),
    .X(net5));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(OUT_1));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(OUT_2));
 sky130_fd_sc_hd__buf_2 fanout8 (.A(net10),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 fanout9 (.A(net10),
    .X(net9));
 sky130_fd_sc_hd__buf_2 fanout10 (.A(wb_clk_i),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 fanout11 (.A(net13),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout12 (.A(net13),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 fanout13 (.A(wb_clk_i),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net12 (.A(net12),
    .X(clknet_0_net12));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net12 (.A(clknet_0_net12),
    .X(clknet_1_0__leaf_net12));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net12 (.A(clknet_0_net12),
    .X(clknet_1_1__leaf_net12));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net8 (.A(net8),
    .X(clknet_0_net8));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net8 (.A(clknet_0_net8),
    .X(clknet_1_0__leaf_net8));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net8 (.A(clknet_0_net8),
    .X(clknet_1_1__leaf_net8));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\count[5] ),
    .X(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(A_PAD));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(B_PAD));
 sky130_fd_sc_hd__diode_2 ANTENNA__1214__B2 (.DIODE(\MUL.PS_R1_inst1.LUT_inst2.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1193__B2 (.DIODE(\MUL.PS_R1_inst1.LUT_inst2.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1044__A1 (.DIODE(\MUL.PS_R1_inst1.LUT_inst2.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0953__A (.DIODE(\MUL.PS_R1_inst1.LUT_inst2.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1166__B2 (.DIODE(\MUL.PS_R1_inst1.LUT_inst3.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__B2 (.DIODE(\MUL.PS_R1_inst1.LUT_inst3.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1025__A1 (.DIODE(\MUL.PS_R1_inst1.LUT_inst3.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0950__A (.DIODE(\MUL.PS_R1_inst1.LUT_inst3.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1138__A1 (.DIODE(\MUL.PS_R1_inst1.LUT_inst4.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1081__B2 (.DIODE(\MUL.PS_R1_inst1.LUT_inst4.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1054__A1 (.DIODE(\MUL.PS_R1_inst1.LUT_inst4.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0946__A (.DIODE(\MUL.PS_R1_inst1.LUT_inst4.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1146__A1 (.DIODE(\MUL.PS_R1_inst1.LUT_inst5.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__A1 (.DIODE(\MUL.PS_R1_inst1.LUT_inst5.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__A1 (.DIODE(\MUL.PS_R1_inst1.LUT_inst5.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0943__A (.DIODE(\MUL.PS_R1_inst1.LUT_inst5.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1090__A1 (.DIODE(\MUL.PS_R1_inst1.LUT_inst6.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1085__A1 (.DIODE(\MUL.PS_R1_inst1.LUT_inst6.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1056__A1 (.DIODE(\MUL.PS_R1_inst1.LUT_inst6.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0940__A (.DIODE(\MUL.PS_R1_inst1.LUT_inst6.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__A1 (.DIODE(\MUL.PS_R1_inst1.LUT_inst8.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1086__A1 (.DIODE(\MUL.PS_R1_inst1.LUT_inst8.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1083__A1 (.DIODE(\MUL.PS_R1_inst1.LUT_inst8.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0932__A (.DIODE(\MUL.PS_R1_inst1.LUT_inst8.I1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__A1 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__A1 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1487__A1 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1486__A1 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1400__B1 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0816__A0 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__S (.DIODE(_0104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1578__S0 (.DIODE(_0104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__S (.DIODE(_0104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1559__B1_N (.DIODE(_0104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1427__B1_N (.DIODE(_0104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__B1 (.DIODE(_0104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1373__B1 (.DIODE(_0104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1335__B1 (.DIODE(_0104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1250__B (.DIODE(_0104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0819__A (.DIODE(_0104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1560__A1 (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1545__S (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1446__B1 (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1345__A1 (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1228__C1 (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__A1 (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__A (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1071__S (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0821__A1 (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0820__A (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1556__A1 (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1555__A1 (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1550__A1_N (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__A1 (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1516__A1 (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1508__B2 (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1504__A1 (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1502__A (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1494__B2 (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0913__B2 (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1556__B2 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__A1 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1524__A1 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__B2 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1512__A1 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__A1_N (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1504__B2 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__A1 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1468__A1 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0917__B2 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__A1 (.DIODE(_0179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__A1_N (.DIODE(_0179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1524__B2 (.DIODE(_0179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__A1 (.DIODE(_0179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1520__A1 (.DIODE(_0179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__B2 (.DIODE(_0179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__B2 (.DIODE(_0179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1458__A1 (.DIODE(_0179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1457__A1 (.DIODE(_0179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0920__A0 (.DIODE(_0179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__B2 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__A1 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1528__A1_N (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__B2 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1477__A1 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1476__A1 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1458__B2 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1432__A1 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1431__A1 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0925__A1 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1540__A1 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__A1_N (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1528__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1477__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__A1 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__A1 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1432__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1403__A1 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1402__A1 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0928__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__B2 (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1466__A1 (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1465__A1_N (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__B2 (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__A1 (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1441__A1 (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1403__B2 (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1391__A1 (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1390__A1 (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0931__B2 (.DIODE(_0187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1348__A1 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1292__B2 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1291__A1 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1172__B2 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__A1 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1130__A1 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1122__B2 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1121__A1 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1087__B2 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0933__A (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__A1 (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__A1_N (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1465__B2 (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__B2 (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1420__A1 (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1419__A1 (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1391__B2 (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1349__A1 (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1306__A1 (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0934__A1 (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__B2 (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1430__A1 (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__A1_N (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1420__B2 (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__A1 (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1393__A1 (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1349__B2 (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1290__A1 (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1289__A1 (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__A0 (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__B2 (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1425__A1 (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1424__A1_N (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__B2 (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1347__A1 (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1346__A1 (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1325__A1 (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1324__A1 (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1290__B2 (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0942__B2 (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1424__B2 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1375__A1 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1374__A1_N (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1346__B2 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1325__B2 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__A1 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1322__A1 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1170__A1 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__A1 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__B2 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1374__B2 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1370__A1 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1369__A1_N (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1331__A1 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1330__A1 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__B2 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1216__B2 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1046__B2 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1025__B2 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0948__A0 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1369__B2 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1288__A1 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1287__A1 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1247__B2 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1246__A1 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1079__B2 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1052__A1 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1051__A1 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1044__B2 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0952__A1 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1340__A1 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1339__A1_N (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1288__B2 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__B2 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1256__A1 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1245__B2 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1225__A1 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__B2 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__A1 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0955__B2 (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1339__B2 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__A1 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1253__A1 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1245__A1 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1225__B2 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1206__A1 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__A1 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__A1 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__B2 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0957__B2 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1580__A1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1273__A1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1268__A1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1263__B (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1261__A2 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1251__B1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1239__B1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1204__B1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__B1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__A0 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0983__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0977__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0976__A (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1308__B1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1267__B (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__B1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1247__B1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1087__B1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1083__B1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1056__B1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1046__B1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1040__B1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__B1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1307__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1256__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1246__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1086__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1055__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1578__A1 (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1259__B1 (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__B1 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1509__A (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1435__A (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1378__A (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1266__B1 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(sel));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout13_A (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout10_A (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0961__A1 (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(wb_rst_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0948__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0934__A0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0924__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0920__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0914__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0904__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__0894__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__0883__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__0880__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__0853__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__0961__S (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1276__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_output7_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1586__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1600__CLK (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__1604__CLK (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout9_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__1615__CLK (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__1633__CLK (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__CLK (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__1638__CLK (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout8_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__1602__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__1614__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__1624__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__1626__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout11_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout12_A (.DIODE(net13));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_617 ();
endmodule

